-- srec2vhdl table generator
-- for input file interrupt_direct.srec

library ieee;
use ieee.std_logic_1164.all;

library work;
use work.processor_common.all;

package processor_common_rom is
    constant rom_contents : rom_type := (
           0 => x"97020000",
           1 => x"93828226",
           2 => x"73905230",
           3 => x"97010020",
           4 => x"9381417f",
           5 => x"17810020",
           6 => x"1301c1fe",
           7 => x"13860188",
           8 => x"93874189",
           9 => x"637af600",
          10 => x"3386c740",
          11 => x"93050000",
          12 => x"13850188",
          13 => x"ef108036",
          14 => x"37050020",
          15 => x"13060500",
          16 => x"93870188",
          17 => x"637cf600",
          18 => x"b7350000",
          19 => x"3386c740",
          20 => x"9385c5fb",
          21 => x"13050500",
          22 => x"ef100032",
          23 => x"ef10006e",
          24 => x"b7050020",
          25 => x"13060000",
          26 => x"93850500",
          27 => x"13055000",
          28 => x"ef104038",
          29 => x"ef108068",
          30 => x"6f00805e",
          31 => x"130101ff",
          32 => x"23261100",
          33 => x"ef008060",
          34 => x"8320c100",
          35 => x"13051000",
          36 => x"13010101",
          37 => x"67800000",
          38 => x"130101fd",
          39 => x"232c4101",
          40 => x"130a0500",
          41 => x"37350000",
          42 => x"130585e0",
          43 => x"23248102",
          44 => x"23229102",
          45 => x"23202103",
          46 => x"232e3101",
          47 => x"83244a08",
          48 => x"23261102",
          49 => x"13044100",
          50 => x"ef00405e",
          51 => x"37390000",
          52 => x"9309c1ff",
          53 => x"93070400",
          54 => x"1309c9bd",
          55 => x"13f7f400",
          56 => x"3307e900",
          57 => x"03470700",
          58 => x"9387f7ff",
          59 => x"93d44400",
          60 => x"2384e700",
          61 => x"e39437ff",
          62 => x"13054100",
          63 => x"23060100",
          64 => x"ef00c05a",
          65 => x"37350000",
          66 => x"1305c5e1",
          67 => x"ef00005a",
          68 => x"03278a08",
          69 => x"9377f700",
          70 => x"b307f900",
          71 => x"83c70700",
          72 => x"1304f4ff",
          73 => x"13574700",
          74 => x"2304f400",
          75 => x"e31434ff",
          76 => x"13054100",
          77 => x"ef008057",
          78 => x"37350000",
          79 => x"130545e5",
          80 => x"ef00c056",
          81 => x"8320c102",
          82 => x"03248102",
          83 => x"83244102",
          84 => x"03290102",
          85 => x"8329c101",
          86 => x"032a8101",
          87 => x"13010103",
          88 => x"67800000",
          89 => x"b70700f0",
          90 => x"03a74708",
          91 => x"1377f7fe",
          92 => x"23a2e708",
          93 => x"03a74700",
          94 => x"13471700",
          95 => x"23a2e700",
          96 => x"67800000",
          97 => x"370700f0",
          98 => x"83274700",
          99 => x"93e70720",
         100 => x"2322f700",
         101 => x"6f000000",
         102 => x"b70700f0",
         103 => x"83a6470f",
         104 => x"03a6070f",
         105 => x"03a7470f",
         106 => x"e31ad7fe",
         107 => x"b7860100",
         108 => x"9305f0ff",
         109 => x"9386066a",
         110 => x"23aeb70e",
         111 => x"b306d600",
         112 => x"23acb70e",
         113 => x"33b6c600",
         114 => x"23acd70e",
         115 => x"3306e600",
         116 => x"23aec70e",
         117 => x"03a74700",
         118 => x"13472700",
         119 => x"23a2e700",
         120 => x"67800000",
         121 => x"b70700f0",
         122 => x"03a74702",
         123 => x"13774700",
         124 => x"630a0700",
         125 => x"03a74700",
         126 => x"13478700",
         127 => x"23a2e700",
         128 => x"83a78702",
         129 => x"67800000",
         130 => x"b70700f0",
         131 => x"03a7470a",
         132 => x"1377f7f0",
         133 => x"23a2e70a",
         134 => x"03a74700",
         135 => x"13474700",
         136 => x"23a2e700",
         137 => x"67800000",
         138 => x"b70700f0",
         139 => x"03a74706",
         140 => x"137777ff",
         141 => x"23a2e706",
         142 => x"03a74700",
         143 => x"13470701",
         144 => x"23a2e700",
         145 => x"67800000",
         146 => x"b70700f0",
         147 => x"03a74704",
         148 => x"137777fe",
         149 => x"23a2e704",
         150 => x"03a74700",
         151 => x"13470702",
         152 => x"23a2e700",
         153 => x"67800000",
         154 => x"6f000000",
         155 => x"13050000",
         156 => x"67800000",
         157 => x"13050000",
         158 => x"67800000",
         159 => x"130101f7",
         160 => x"23221100",
         161 => x"23242100",
         162 => x"23263100",
         163 => x"23284100",
         164 => x"232a5100",
         165 => x"232c6100",
         166 => x"232e7100",
         167 => x"23208102",
         168 => x"23229102",
         169 => x"2324a102",
         170 => x"2326b102",
         171 => x"2328c102",
         172 => x"232ad102",
         173 => x"232ce102",
         174 => x"232ef102",
         175 => x"23200105",
         176 => x"23221105",
         177 => x"23242105",
         178 => x"23263105",
         179 => x"23284105",
         180 => x"232a5105",
         181 => x"232c6105",
         182 => x"232e7105",
         183 => x"23208107",
         184 => x"23229107",
         185 => x"2324a107",
         186 => x"2326b107",
         187 => x"2328c107",
         188 => x"232ad107",
         189 => x"232ce107",
         190 => x"232ef107",
         191 => x"f3222034",
         192 => x"23205108",
         193 => x"f3221034",
         194 => x"23225108",
         195 => x"83a20200",
         196 => x"23245108",
         197 => x"f3223034",
         198 => x"23265108",
         199 => x"f3272034",
         200 => x"37070080",
         201 => x"93067700",
         202 => x"6386d70e",
         203 => x"9306b000",
         204 => x"63fef602",
         205 => x"934607ff",
         206 => x"b386d700",
         207 => x"13065000",
         208 => x"636ad602",
         209 => x"1347f7fe",
         210 => x"b387e700",
         211 => x"13074000",
         212 => x"636af714",
         213 => x"37370000",
         214 => x"93972700",
         215 => x"130707bf",
         216 => x"b387e700",
         217 => x"83a70700",
         218 => x"67800700",
         219 => x"13071000",
         220 => x"6364f708",
         221 => x"03258102",
         222 => x"832fc107",
         223 => x"032f8107",
         224 => x"832e4107",
         225 => x"032e0107",
         226 => x"832dc106",
         227 => x"032d8106",
         228 => x"832c4106",
         229 => x"032c0106",
         230 => x"832bc105",
         231 => x"032b8105",
         232 => x"832a4105",
         233 => x"032a0105",
         234 => x"8329c104",
         235 => x"03298104",
         236 => x"83284104",
         237 => x"03280104",
         238 => x"8327c103",
         239 => x"03278103",
         240 => x"83264103",
         241 => x"03260103",
         242 => x"8325c102",
         243 => x"83244102",
         244 => x"03240102",
         245 => x"8323c101",
         246 => x"03238101",
         247 => x"83224101",
         248 => x"03220101",
         249 => x"8321c100",
         250 => x"03218100",
         251 => x"83204100",
         252 => x"13010109",
         253 => x"73002030",
         254 => x"e3eef6f6",
         255 => x"37370000",
         256 => x"93972700",
         257 => x"130747c0",
         258 => x"b387e700",
         259 => x"83a70700",
         260 => x"67800700",
         261 => x"eff05fd8",
         262 => x"03258102",
         263 => x"6ff0dff5",
         264 => x"eff09fde",
         265 => x"03258102",
         266 => x"6ff01ff5",
         267 => x"eff0dfdf",
         268 => x"03258102",
         269 => x"6ff05ff4",
         270 => x"eff01fe1",
         271 => x"03258102",
         272 => x"6ff09ff3",
         273 => x"eff01fd2",
         274 => x"03258102",
         275 => x"6ff0dff2",
         276 => x"eff05fd9",
         277 => x"03258102",
         278 => x"6ff01ff2",
         279 => x"9307600d",
         280 => x"6384f806",
         281 => x"9307900a",
         282 => x"6388f818",
         283 => x"63ca170f",
         284 => x"938878fc",
         285 => x"93074002",
         286 => x"63ec1703",
         287 => x"b7370000",
         288 => x"938747c3",
         289 => x"93982800",
         290 => x"b388f800",
         291 => x"83a70800",
         292 => x"67800700",
         293 => x"13050100",
         294 => x"eff01fc0",
         295 => x"03258102",
         296 => x"6ff09fed",
         297 => x"eff01fce",
         298 => x"03258102",
         299 => x"6ff0dfec",
         300 => x"ef104024",
         301 => x"93078005",
         302 => x"2320f500",
         303 => x"9307f0ff",
         304 => x"13850700",
         305 => x"6ff05feb",
         306 => x"63120510",
         307 => x"13858189",
         308 => x"13050500",
         309 => x"6ff05fea",
         310 => x"b7270000",
         311 => x"23a2f500",
         312 => x"93070000",
         313 => x"13850700",
         314 => x"6ff01fe9",
         315 => x"93070000",
         316 => x"13850700",
         317 => x"6ff05fe8",
         318 => x"ef10c01f",
         319 => x"93079000",
         320 => x"2320f500",
         321 => x"9307f0ff",
         322 => x"13850700",
         323 => x"6ff0dfe6",
         324 => x"13090600",
         325 => x"13840500",
         326 => x"635cc000",
         327 => x"b384c500",
         328 => x"03450400",
         329 => x"13041400",
         330 => x"eff05fb5",
         331 => x"e39a84fe",
         332 => x"13050900",
         333 => x"6ff05fe4",
         334 => x"13090600",
         335 => x"13840500",
         336 => x"e358c0fe",
         337 => x"b384c500",
         338 => x"eff01fb3",
         339 => x"2300a400",
         340 => x"13041400",
         341 => x"e31a94fe",
         342 => x"13050900",
         343 => x"6ff0dfe1",
         344 => x"938808c0",
         345 => x"9307f000",
         346 => x"e3e417f5",
         347 => x"b7370000",
         348 => x"938787cc",
         349 => x"93982800",
         350 => x"b388f800",
         351 => x"83a70800",
         352 => x"67800700",
         353 => x"ef100017",
         354 => x"9307d000",
         355 => x"2320f500",
         356 => x"9307f0ff",
         357 => x"13850700",
         358 => x"6ff01fde",
         359 => x"ef108015",
         360 => x"93072000",
         361 => x"2320f500",
         362 => x"9307f0ff",
         363 => x"13850700",
         364 => x"6ff09fdc",
         365 => x"ef100014",
         366 => x"9307f001",
         367 => x"2320f500",
         368 => x"9307f0ff",
         369 => x"13850700",
         370 => x"6ff01fdb",
         371 => x"b7870020",
         372 => x"93870700",
         373 => x"13070040",
         374 => x"b387e740",
         375 => x"e36af5ee",
         376 => x"ef104011",
         377 => x"9307c000",
         378 => x"2320f500",
         379 => x"1305f0ff",
         380 => x"13050500",
         381 => x"6ff05fd8",
         382 => x"13090000",
         383 => x"93040500",
         384 => x"13040900",
         385 => x"93090900",
         386 => x"93070900",
         387 => x"732410c8",
         388 => x"f32910c0",
         389 => x"f32710c8",
         390 => x"e31af4fe",
         391 => x"37460f00",
         392 => x"13060624",
         393 => x"93060000",
         394 => x"13850900",
         395 => x"93050400",
         396 => x"ef005016",
         397 => x"37460f00",
         398 => x"23a4a400",
         399 => x"13060624",
         400 => x"93060000",
         401 => x"13850900",
         402 => x"93050400",
         403 => x"ef008051",
         404 => x"23a0a400",
         405 => x"23a2b400",
         406 => x"13050900",
         407 => x"6ff0dfd1",
         408 => x"370700f0",
         409 => x"83274702",
         410 => x"93f74700",
         411 => x"e38c07fe",
         412 => x"03258702",
         413 => x"1375f50f",
         414 => x"67800000",
         415 => x"b70700f0",
         416 => x"23a6a702",
         417 => x"23a0b702",
         418 => x"67800000",
         419 => x"1375f50f",
         420 => x"b70700f0",
         421 => x"370700f0",
         422 => x"23a4a702",
         423 => x"83274702",
         424 => x"93f70701",
         425 => x"e38c07fe",
         426 => x"67800000",
         427 => x"630e0502",
         428 => x"130101ff",
         429 => x"23248100",
         430 => x"23261100",
         431 => x"13040500",
         432 => x"03450500",
         433 => x"630a0500",
         434 => x"13041400",
         435 => x"eff01ffc",
         436 => x"03450400",
         437 => x"e31a05fe",
         438 => x"8320c100",
         439 => x"03248100",
         440 => x"13010101",
         441 => x"67800000",
         442 => x"67800000",
         443 => x"13030500",
         444 => x"138e0500",
         445 => x"93080000",
         446 => x"63dc0500",
         447 => x"b337a000",
         448 => x"330eb040",
         449 => x"330efe40",
         450 => x"3303a040",
         451 => x"9308f0ff",
         452 => x"63dc0600",
         453 => x"b337c000",
         454 => x"b306d040",
         455 => x"93c8f8ff",
         456 => x"b386f640",
         457 => x"3306c040",
         458 => x"13070600",
         459 => x"13080300",
         460 => x"93070e00",
         461 => x"639c0628",
         462 => x"b7350000",
         463 => x"938585d0",
         464 => x"6376ce0e",
         465 => x"b7060100",
         466 => x"6378d60c",
         467 => x"93360610",
         468 => x"93c61600",
         469 => x"93963600",
         470 => x"3355d600",
         471 => x"b385a500",
         472 => x"83c50500",
         473 => x"13050002",
         474 => x"b386d500",
         475 => x"b305d540",
         476 => x"630cd500",
         477 => x"b317be00",
         478 => x"b356d300",
         479 => x"3317b600",
         480 => x"b3e7f600",
         481 => x"3318b300",
         482 => x"93550701",
         483 => x"33deb702",
         484 => x"13160701",
         485 => x"13560601",
         486 => x"b3f7b702",
         487 => x"13050e00",
         488 => x"3303c603",
         489 => x"93960701",
         490 => x"93570801",
         491 => x"b3e7d700",
         492 => x"63fe6700",
         493 => x"b307f700",
         494 => x"1305feff",
         495 => x"63e8e700",
         496 => x"63f66700",
         497 => x"1305eeff",
         498 => x"b387e700",
         499 => x"b3876740",
         500 => x"33d3b702",
         501 => x"13180801",
         502 => x"13580801",
         503 => x"b3f7b702",
         504 => x"b3066602",
         505 => x"93970701",
         506 => x"3368f800",
         507 => x"93070300",
         508 => x"637cd800",
         509 => x"33080701",
         510 => x"9307f3ff",
         511 => x"6366e800",
         512 => x"6374d800",
         513 => x"9307e3ff",
         514 => x"13150501",
         515 => x"3365f500",
         516 => x"93050000",
         517 => x"6f00000e",
         518 => x"37050001",
         519 => x"93060001",
         520 => x"e36ca6f2",
         521 => x"93068001",
         522 => x"6ff01ff3",
         523 => x"93060000",
         524 => x"630c0600",
         525 => x"b7070100",
         526 => x"637af60c",
         527 => x"93360610",
         528 => x"93c61600",
         529 => x"93963600",
         530 => x"b357d600",
         531 => x"b385f500",
         532 => x"83c70500",
         533 => x"b387d700",
         534 => x"93060002",
         535 => x"b385f640",
         536 => x"6390f60c",
         537 => x"b307ce40",
         538 => x"93051000",
         539 => x"13530701",
         540 => x"b3de6702",
         541 => x"13160701",
         542 => x"13560601",
         543 => x"93560801",
         544 => x"b3f76702",
         545 => x"13850e00",
         546 => x"330ed603",
         547 => x"93970701",
         548 => x"b3e7f600",
         549 => x"63fec701",
         550 => x"b307f700",
         551 => x"1385feff",
         552 => x"63e8e700",
         553 => x"63f6c701",
         554 => x"1385eeff",
         555 => x"b387e700",
         556 => x"b387c741",
         557 => x"33de6702",
         558 => x"13180801",
         559 => x"13580801",
         560 => x"b3f76702",
         561 => x"b306c603",
         562 => x"93970701",
         563 => x"3368f800",
         564 => x"93070e00",
         565 => x"637cd800",
         566 => x"33080701",
         567 => x"9307feff",
         568 => x"6366e800",
         569 => x"6374d800",
         570 => x"9307eeff",
         571 => x"13150501",
         572 => x"3365f500",
         573 => x"638a0800",
         574 => x"b337a000",
         575 => x"b305b040",
         576 => x"b385f540",
         577 => x"3305a040",
         578 => x"67800000",
         579 => x"b7070001",
         580 => x"93060001",
         581 => x"e36af6f2",
         582 => x"93068001",
         583 => x"6ff0dff2",
         584 => x"3317b600",
         585 => x"b356fe00",
         586 => x"13550701",
         587 => x"331ebe00",
         588 => x"b357f300",
         589 => x"b3e7c701",
         590 => x"33dea602",
         591 => x"13160701",
         592 => x"13560601",
         593 => x"3318b300",
         594 => x"b3f6a602",
         595 => x"3303c603",
         596 => x"93950601",
         597 => x"93d60701",
         598 => x"b3e6b600",
         599 => x"93050e00",
         600 => x"63fe6600",
         601 => x"b306d700",
         602 => x"9305feff",
         603 => x"63e8e600",
         604 => x"63f66600",
         605 => x"9305eeff",
         606 => x"b386e600",
         607 => x"b3866640",
         608 => x"33d3a602",
         609 => x"93970701",
         610 => x"93d70701",
         611 => x"b3f6a602",
         612 => x"33066602",
         613 => x"93960601",
         614 => x"b3e7d700",
         615 => x"93060300",
         616 => x"63fec700",
         617 => x"b307f700",
         618 => x"9306f3ff",
         619 => x"63e8e700",
         620 => x"63f6c700",
         621 => x"9306e3ff",
         622 => x"b387e700",
         623 => x"93950501",
         624 => x"b387c740",
         625 => x"b3e5d500",
         626 => x"6ff05fea",
         627 => x"6366de18",
         628 => x"b7070100",
         629 => x"63f4f604",
         630 => x"13b70610",
         631 => x"13471700",
         632 => x"13173700",
         633 => x"b7370000",
         634 => x"b3d5e600",
         635 => x"938787d0",
         636 => x"b387b700",
         637 => x"83c70700",
         638 => x"b387e700",
         639 => x"13070002",
         640 => x"b305f740",
         641 => x"6316f702",
         642 => x"13051000",
         643 => x"e3e4c6ef",
         644 => x"3335c300",
         645 => x"13451500",
         646 => x"6ff0dfed",
         647 => x"b7070001",
         648 => x"13070001",
         649 => x"e3e0f6fc",
         650 => x"13078001",
         651 => x"6ff09ffb",
         652 => x"3357f600",
         653 => x"b396b600",
         654 => x"b366d700",
         655 => x"3357fe00",
         656 => x"331ebe00",
         657 => x"b357f300",
         658 => x"b3e7c701",
         659 => x"13de0601",
         660 => x"335fc703",
         661 => x"13980601",
         662 => x"13580801",
         663 => x"3316b600",
         664 => x"3377c703",
         665 => x"b30ee803",
         666 => x"13150701",
         667 => x"13d70701",
         668 => x"3367a700",
         669 => x"13050f00",
         670 => x"637ed701",
         671 => x"3387e600",
         672 => x"1305ffff",
         673 => x"6368d700",
         674 => x"6376d701",
         675 => x"1305efff",
         676 => x"3307d700",
         677 => x"3307d741",
         678 => x"b35ec703",
         679 => x"93970701",
         680 => x"93d70701",
         681 => x"3377c703",
         682 => x"3308d803",
         683 => x"13170701",
         684 => x"b3e7e700",
         685 => x"13870e00",
         686 => x"63fe0701",
         687 => x"b387f600",
         688 => x"1387feff",
         689 => x"63e8d700",
         690 => x"63f60701",
         691 => x"1387eeff",
         692 => x"b387d700",
         693 => x"13150501",
         694 => x"b70e0100",
         695 => x"3365e500",
         696 => x"9386feff",
         697 => x"3377d500",
         698 => x"b3870741",
         699 => x"b376d600",
         700 => x"13580501",
         701 => x"13560601",
         702 => x"330ed702",
         703 => x"b306d802",
         704 => x"3307c702",
         705 => x"3308c802",
         706 => x"3306d700",
         707 => x"13570e01",
         708 => x"3307c700",
         709 => x"6374d700",
         710 => x"3308d801",
         711 => x"93560701",
         712 => x"b3860601",
         713 => x"63e6d702",
         714 => x"e394d7ce",
         715 => x"b7070100",
         716 => x"9387f7ff",
         717 => x"3377f700",
         718 => x"13170701",
         719 => x"337efe00",
         720 => x"3313b300",
         721 => x"3307c701",
         722 => x"93050000",
         723 => x"e374e3da",
         724 => x"1305f5ff",
         725 => x"6ff0dfcb",
         726 => x"93050000",
         727 => x"13050000",
         728 => x"6ff05fd9",
         729 => x"93080500",
         730 => x"13830500",
         731 => x"13070600",
         732 => x"13080500",
         733 => x"93870500",
         734 => x"63920628",
         735 => x"b7350000",
         736 => x"938585d0",
         737 => x"6376c30e",
         738 => x"b7060100",
         739 => x"6378d60c",
         740 => x"93360610",
         741 => x"93c61600",
         742 => x"93963600",
         743 => x"3355d600",
         744 => x"b385a500",
         745 => x"83c50500",
         746 => x"13050002",
         747 => x"b386d500",
         748 => x"b305d540",
         749 => x"630cd500",
         750 => x"b317b300",
         751 => x"b3d6d800",
         752 => x"3317b600",
         753 => x"b3e7f600",
         754 => x"3398b800",
         755 => x"93550701",
         756 => x"33d3b702",
         757 => x"13160701",
         758 => x"13560601",
         759 => x"b3f7b702",
         760 => x"13050300",
         761 => x"b3086602",
         762 => x"93960701",
         763 => x"93570801",
         764 => x"b3e7d700",
         765 => x"63fe1701",
         766 => x"b307f700",
         767 => x"1305f3ff",
         768 => x"63e8e700",
         769 => x"63f61701",
         770 => x"1305e3ff",
         771 => x"b387e700",
         772 => x"b3871741",
         773 => x"b3d8b702",
         774 => x"13180801",
         775 => x"13580801",
         776 => x"b3f7b702",
         777 => x"b3061603",
         778 => x"93970701",
         779 => x"3368f800",
         780 => x"93870800",
         781 => x"637cd800",
         782 => x"33080701",
         783 => x"9387f8ff",
         784 => x"6366e800",
         785 => x"6374d800",
         786 => x"9387e8ff",
         787 => x"13150501",
         788 => x"3365f500",
         789 => x"93050000",
         790 => x"67800000",
         791 => x"37050001",
         792 => x"93060001",
         793 => x"e36ca6f2",
         794 => x"93068001",
         795 => x"6ff01ff3",
         796 => x"93060000",
         797 => x"630c0600",
         798 => x"b7070100",
         799 => x"6370f60c",
         800 => x"93360610",
         801 => x"93c61600",
         802 => x"93963600",
         803 => x"b357d600",
         804 => x"b385f500",
         805 => x"83c70500",
         806 => x"b387d700",
         807 => x"93060002",
         808 => x"b385f640",
         809 => x"6396f60a",
         810 => x"b307c340",
         811 => x"93051000",
         812 => x"93580701",
         813 => x"33de1703",
         814 => x"13160701",
         815 => x"13560601",
         816 => x"93560801",
         817 => x"b3f71703",
         818 => x"13050e00",
         819 => x"3303c603",
         820 => x"93970701",
         821 => x"b3e7f600",
         822 => x"63fe6700",
         823 => x"b307f700",
         824 => x"1305feff",
         825 => x"63e8e700",
         826 => x"63f66700",
         827 => x"1305eeff",
         828 => x"b387e700",
         829 => x"b3876740",
         830 => x"33d31703",
         831 => x"13180801",
         832 => x"13580801",
         833 => x"b3f71703",
         834 => x"b3066602",
         835 => x"93970701",
         836 => x"3368f800",
         837 => x"93070300",
         838 => x"637cd800",
         839 => x"33080701",
         840 => x"9307f3ff",
         841 => x"6366e800",
         842 => x"6374d800",
         843 => x"9307e3ff",
         844 => x"13150501",
         845 => x"3365f500",
         846 => x"67800000",
         847 => x"b7070001",
         848 => x"93060001",
         849 => x"e364f6f4",
         850 => x"93068001",
         851 => x"6ff01ff4",
         852 => x"3317b600",
         853 => x"b356f300",
         854 => x"13550701",
         855 => x"3313b300",
         856 => x"b3d7f800",
         857 => x"b3e76700",
         858 => x"33d3a602",
         859 => x"13160701",
         860 => x"13560601",
         861 => x"3398b800",
         862 => x"b3f6a602",
         863 => x"b3086602",
         864 => x"93950601",
         865 => x"93d60701",
         866 => x"b3e6b600",
         867 => x"93050300",
         868 => x"63fe1601",
         869 => x"b306d700",
         870 => x"9305f3ff",
         871 => x"63e8e600",
         872 => x"63f61601",
         873 => x"9305e3ff",
         874 => x"b386e600",
         875 => x"b3861641",
         876 => x"b3d8a602",
         877 => x"93970701",
         878 => x"93d70701",
         879 => x"b3f6a602",
         880 => x"33061603",
         881 => x"93960601",
         882 => x"b3e7d700",
         883 => x"93860800",
         884 => x"63fec700",
         885 => x"b307f700",
         886 => x"9386f8ff",
         887 => x"63e8e700",
         888 => x"63f6c700",
         889 => x"9386e8ff",
         890 => x"b387e700",
         891 => x"93950501",
         892 => x"b387c740",
         893 => x"b3e5d500",
         894 => x"6ff09feb",
         895 => x"63e6d518",
         896 => x"b7070100",
         897 => x"63f4f604",
         898 => x"13b70610",
         899 => x"13471700",
         900 => x"13173700",
         901 => x"b7370000",
         902 => x"b3d5e600",
         903 => x"938787d0",
         904 => x"b387b700",
         905 => x"83c70700",
         906 => x"b387e700",
         907 => x"13070002",
         908 => x"b305f740",
         909 => x"6316f702",
         910 => x"13051000",
         911 => x"e3ee66e0",
         912 => x"33b5c800",
         913 => x"13451500",
         914 => x"67800000",
         915 => x"b7070001",
         916 => x"13070001",
         917 => x"e3e0f6fc",
         918 => x"13078001",
         919 => x"6ff09ffb",
         920 => x"3357f600",
         921 => x"b396b600",
         922 => x"b366d700",
         923 => x"3357f300",
         924 => x"3313b300",
         925 => x"b3d7f800",
         926 => x"b3e76700",
         927 => x"13d30601",
         928 => x"b35e6702",
         929 => x"13980601",
         930 => x"13580801",
         931 => x"3316b600",
         932 => x"33776702",
         933 => x"330ed803",
         934 => x"13150701",
         935 => x"13d70701",
         936 => x"3367a700",
         937 => x"13850e00",
         938 => x"637ec701",
         939 => x"3387e600",
         940 => x"1385feff",
         941 => x"6368d700",
         942 => x"6376c701",
         943 => x"1385eeff",
         944 => x"3307d700",
         945 => x"3307c741",
         946 => x"335e6702",
         947 => x"93970701",
         948 => x"93d70701",
         949 => x"33776702",
         950 => x"3308c803",
         951 => x"13170701",
         952 => x"b3e7e700",
         953 => x"13070e00",
         954 => x"63fe0701",
         955 => x"b387f600",
         956 => x"1307feff",
         957 => x"63e8d700",
         958 => x"63f60701",
         959 => x"1307eeff",
         960 => x"b387d700",
         961 => x"13150501",
         962 => x"370e0100",
         963 => x"3365e500",
         964 => x"9306feff",
         965 => x"3377d500",
         966 => x"b3870741",
         967 => x"b376d600",
         968 => x"13580501",
         969 => x"13560601",
         970 => x"3303d702",
         971 => x"b306d802",
         972 => x"3307c702",
         973 => x"3308c802",
         974 => x"3306d700",
         975 => x"13570301",
         976 => x"3307c700",
         977 => x"6374d700",
         978 => x"3308c801",
         979 => x"93560701",
         980 => x"b3860601",
         981 => x"63e6d702",
         982 => x"e39ed7ce",
         983 => x"b7070100",
         984 => x"9387f7ff",
         985 => x"3377f700",
         986 => x"13170701",
         987 => x"3373f300",
         988 => x"b398b800",
         989 => x"33076700",
         990 => x"93050000",
         991 => x"e3fee8cc",
         992 => x"1305f5ff",
         993 => x"6ff01fcd",
         994 => x"93050000",
         995 => x"13050000",
         996 => x"67800000",
         997 => x"13080600",
         998 => x"93070500",
         999 => x"13870500",
        1000 => x"63960620",
        1001 => x"b7380000",
        1002 => x"938888d0",
        1003 => x"63fcc50c",
        1004 => x"b7060100",
        1005 => x"637ed60a",
        1006 => x"93360610",
        1007 => x"93c61600",
        1008 => x"93963600",
        1009 => x"3353d600",
        1010 => x"b3886800",
        1011 => x"83c80800",
        1012 => x"13030002",
        1013 => x"b386d800",
        1014 => x"b308d340",
        1015 => x"630cd300",
        1016 => x"33971501",
        1017 => x"b356d500",
        1018 => x"33181601",
        1019 => x"33e7e600",
        1020 => x"b3171501",
        1021 => x"13560801",
        1022 => x"b356c702",
        1023 => x"13150801",
        1024 => x"13550501",
        1025 => x"3377c702",
        1026 => x"b386a602",
        1027 => x"93150701",
        1028 => x"13d70701",
        1029 => x"3367b700",
        1030 => x"637ad700",
        1031 => x"3307e800",
        1032 => x"63660701",
        1033 => x"6374d700",
        1034 => x"33070701",
        1035 => x"3307d740",
        1036 => x"b356c702",
        1037 => x"3377c702",
        1038 => x"b386a602",
        1039 => x"93970701",
        1040 => x"13170701",
        1041 => x"93d70701",
        1042 => x"b3e7e700",
        1043 => x"63fad700",
        1044 => x"b307f800",
        1045 => x"63e60701",
        1046 => x"63f4d700",
        1047 => x"b3870701",
        1048 => x"b387d740",
        1049 => x"33d51701",
        1050 => x"93050000",
        1051 => x"67800000",
        1052 => x"37030001",
        1053 => x"93060001",
        1054 => x"e36666f4",
        1055 => x"93068001",
        1056 => x"6ff05ff4",
        1057 => x"93060000",
        1058 => x"630c0600",
        1059 => x"37070100",
        1060 => x"637ee606",
        1061 => x"93360610",
        1062 => x"93c61600",
        1063 => x"93963600",
        1064 => x"3357d600",
        1065 => x"b388e800",
        1066 => x"03c70800",
        1067 => x"3307d700",
        1068 => x"93060002",
        1069 => x"b388e640",
        1070 => x"6394e606",
        1071 => x"3387c540",
        1072 => x"93550801",
        1073 => x"3356b702",
        1074 => x"13150801",
        1075 => x"13550501",
        1076 => x"93d60701",
        1077 => x"3377b702",
        1078 => x"3306a602",
        1079 => x"13170701",
        1080 => x"33e7e600",
        1081 => x"637ac700",
        1082 => x"3307e800",
        1083 => x"63660701",
        1084 => x"6374c700",
        1085 => x"33070701",
        1086 => x"3307c740",
        1087 => x"b356b702",
        1088 => x"3377b702",
        1089 => x"b386a602",
        1090 => x"6ff05ff3",
        1091 => x"37070001",
        1092 => x"93060001",
        1093 => x"e366e6f8",
        1094 => x"93068001",
        1095 => x"6ff05ff8",
        1096 => x"33181601",
        1097 => x"b3d6e500",
        1098 => x"b3171501",
        1099 => x"b3951501",
        1100 => x"3357e500",
        1101 => x"13550801",
        1102 => x"3367b700",
        1103 => x"b3d5a602",
        1104 => x"13130801",
        1105 => x"13530301",
        1106 => x"b3f6a602",
        1107 => x"b3856502",
        1108 => x"13960601",
        1109 => x"93560701",
        1110 => x"b3e6c600",
        1111 => x"63fab600",
        1112 => x"b306d800",
        1113 => x"63e60601",
        1114 => x"63f4b600",
        1115 => x"b3860601",
        1116 => x"b386b640",
        1117 => x"33d6a602",
        1118 => x"13170701",
        1119 => x"13570701",
        1120 => x"b3f6a602",
        1121 => x"33066602",
        1122 => x"93960601",
        1123 => x"3367d700",
        1124 => x"637ac700",
        1125 => x"3307e800",
        1126 => x"63660701",
        1127 => x"6374c700",
        1128 => x"33070701",
        1129 => x"3307c740",
        1130 => x"6ff09ff1",
        1131 => x"63e4d51c",
        1132 => x"37080100",
        1133 => x"63fe0605",
        1134 => x"13b80610",
        1135 => x"13481800",
        1136 => x"13183800",
        1137 => x"b7380000",
        1138 => x"33d30601",
        1139 => x"938888d0",
        1140 => x"b3886800",
        1141 => x"83c80800",
        1142 => x"13030002",
        1143 => x"b3880801",
        1144 => x"33081341",
        1145 => x"63101305",
        1146 => x"63e4b600",
        1147 => x"636cc500",
        1148 => x"3306c540",
        1149 => x"b386d540",
        1150 => x"3337c500",
        1151 => x"93070600",
        1152 => x"3387e640",
        1153 => x"13850700",
        1154 => x"93050700",
        1155 => x"67800000",
        1156 => x"b7080001",
        1157 => x"13080001",
        1158 => x"e3e616fb",
        1159 => x"13088001",
        1160 => x"6ff05ffa",
        1161 => x"b3571601",
        1162 => x"b3960601",
        1163 => x"b3e6d700",
        1164 => x"33d71501",
        1165 => x"13de0601",
        1166 => x"335fc703",
        1167 => x"13930601",
        1168 => x"13530301",
        1169 => x"b3970501",
        1170 => x"b3551501",
        1171 => x"b3e5f500",
        1172 => x"93d70501",
        1173 => x"33160601",
        1174 => x"33150501",
        1175 => x"3377c703",
        1176 => x"b30ee303",
        1177 => x"13170701",
        1178 => x"b3e7e700",
        1179 => x"13070f00",
        1180 => x"63fed701",
        1181 => x"b387f600",
        1182 => x"1307ffff",
        1183 => x"63e8d700",
        1184 => x"63f6d701",
        1185 => x"1307efff",
        1186 => x"b387d700",
        1187 => x"b387d741",
        1188 => x"b3dec703",
        1189 => x"93950501",
        1190 => x"93d50501",
        1191 => x"b3f7c703",
        1192 => x"138e0e00",
        1193 => x"3303d303",
        1194 => x"93970701",
        1195 => x"b3e5f500",
        1196 => x"63fe6500",
        1197 => x"b385b600",
        1198 => x"138efeff",
        1199 => x"63e8d500",
        1200 => x"63f66500",
        1201 => x"138eeeff",
        1202 => x"b385d500",
        1203 => x"93170701",
        1204 => x"370f0100",
        1205 => x"b3e7c701",
        1206 => x"b3856540",
        1207 => x"1303ffff",
        1208 => x"33f76700",
        1209 => x"135e0601",
        1210 => x"93d70701",
        1211 => x"33736600",
        1212 => x"b30e6702",
        1213 => x"33836702",
        1214 => x"3307c703",
        1215 => x"b387c703",
        1216 => x"330e6700",
        1217 => x"13d70e01",
        1218 => x"3307c701",
        1219 => x"63746700",
        1220 => x"b387e701",
        1221 => x"13530701",
        1222 => x"b307f300",
        1223 => x"37030100",
        1224 => x"1303f3ff",
        1225 => x"33776700",
        1226 => x"13170701",
        1227 => x"b3fe6e00",
        1228 => x"3307d701",
        1229 => x"63e6f500",
        1230 => x"639ef500",
        1231 => x"637ce500",
        1232 => x"3306c740",
        1233 => x"3333c700",
        1234 => x"b306d300",
        1235 => x"13070600",
        1236 => x"b387d740",
        1237 => x"3307e540",
        1238 => x"3335e500",
        1239 => x"b385f540",
        1240 => x"b385a540",
        1241 => x"b3981501",
        1242 => x"33570701",
        1243 => x"33e5e800",
        1244 => x"b3d50501",
        1245 => x"67800000",
        1246 => x"13030500",
        1247 => x"630e0600",
        1248 => x"83830500",
        1249 => x"23007300",
        1250 => x"1306f6ff",
        1251 => x"13031300",
        1252 => x"93851500",
        1253 => x"e31606fe",
        1254 => x"67800000",
        1255 => x"13030500",
        1256 => x"630a0600",
        1257 => x"2300b300",
        1258 => x"1306f6ff",
        1259 => x"13031300",
        1260 => x"e31a06fe",
        1261 => x"67800000",
        1262 => x"630c0602",
        1263 => x"13030500",
        1264 => x"93061000",
        1265 => x"636ab500",
        1266 => x"9306f0ff",
        1267 => x"1307f6ff",
        1268 => x"3303e300",
        1269 => x"b385e500",
        1270 => x"83830500",
        1271 => x"23007300",
        1272 => x"1306f6ff",
        1273 => x"3303d300",
        1274 => x"b385d500",
        1275 => x"e31606fe",
        1276 => x"67800000",
        1277 => x"130101f9",
        1278 => x"23248106",
        1279 => x"23229106",
        1280 => x"23261106",
        1281 => x"23202107",
        1282 => x"232e3105",
        1283 => x"232c4105",
        1284 => x"232a5105",
        1285 => x"23286105",
        1286 => x"23267105",
        1287 => x"23248105",
        1288 => x"23229105",
        1289 => x"2320a105",
        1290 => x"93040500",
        1291 => x"13840500",
        1292 => x"232c0100",
        1293 => x"232e0100",
        1294 => x"23200102",
        1295 => x"23220102",
        1296 => x"23240102",
        1297 => x"23260102",
        1298 => x"23280102",
        1299 => x"232a0102",
        1300 => x"232c0102",
        1301 => x"232e0102",
        1302 => x"97f2ffff",
        1303 => x"938242e2",
        1304 => x"73905230",
        1305 => x"93050004",
        1306 => x"1305101b",
        1307 => x"eff00fa1",
        1308 => x"37877d01",
        1309 => x"b70700f0",
        1310 => x"1307f783",
        1311 => x"23a6e708",
        1312 => x"93061001",
        1313 => x"37170000",
        1314 => x"23a0d708",
        1315 => x"13077738",
        1316 => x"23a8e70a",
        1317 => x"37270000",
        1318 => x"1307f770",
        1319 => x"23a6e70a",
        1320 => x"23a0d70a",
        1321 => x"13078070",
        1322 => x"23a0e706",
        1323 => x"3707f900",
        1324 => x"13078700",
        1325 => x"23a0e704",
        1326 => x"93020008",
        1327 => x"73904230",
        1328 => x"b7220000",
        1329 => x"93828280",
        1330 => x"73900230",
        1331 => x"b7390000",
        1332 => x"138549e5",
        1333 => x"eff08f9d",
        1334 => x"63549002",
        1335 => x"1389f4ff",
        1336 => x"9304f0ff",
        1337 => x"03250400",
        1338 => x"1309f9ff",
        1339 => x"13044400",
        1340 => x"eff0cf9b",
        1341 => x"138549e5",
        1342 => x"eff04f9b",
        1343 => x"e31499fe",
        1344 => x"37350000",
        1345 => x"b7faeeee",
        1346 => x"130585e2",
        1347 => x"b7090010",
        1348 => x"37140000",
        1349 => x"1389faee",
        1350 => x"eff04f99",
        1351 => x"373b0000",
        1352 => x"9389f9ff",
        1353 => x"938aeaee",
        1354 => x"130404e1",
        1355 => x"93040000",
        1356 => x"b71b0000",
        1357 => x"938b0b2c",
        1358 => x"130af000",
        1359 => x"93050000",
        1360 => x"13058100",
        1361 => x"ef008036",
        1362 => x"938bfbff",
        1363 => x"630a0502",
        1364 => x"e3960bfe",
        1365 => x"73001000",
        1366 => x"b70700f0",
        1367 => x"9306f00f",
        1368 => x"23a4d706",
        1369 => x"03a70704",
        1370 => x"93860704",
        1371 => x"13670730",
        1372 => x"23a0e704",
        1373 => x"93070009",
        1374 => x"23a4f600",
        1375 => x"6ff05ffb",
        1376 => x"032c8100",
        1377 => x"8325c100",
        1378 => x"13060400",
        1379 => x"9357cc01",
        1380 => x"13974500",
        1381 => x"b367f700",
        1382 => x"b3f73701",
        1383 => x"33773c01",
        1384 => x"13d5f541",
        1385 => x"13d88501",
        1386 => x"3307f700",
        1387 => x"33070701",
        1388 => x"9377d500",
        1389 => x"3307f700",
        1390 => x"33774703",
        1391 => x"937725ff",
        1392 => x"93860400",
        1393 => x"13050c00",
        1394 => x"3307f700",
        1395 => x"b307ec40",
        1396 => x"1357f741",
        1397 => x"3338fc00",
        1398 => x"3387e540",
        1399 => x"33070741",
        1400 => x"b3885703",
        1401 => x"33072703",
        1402 => x"33b82703",
        1403 => x"33071701",
        1404 => x"b3872703",
        1405 => x"33070701",
        1406 => x"1358f741",
        1407 => x"13783800",
        1408 => x"b307f800",
        1409 => x"33b80701",
        1410 => x"3307e800",
        1411 => x"1318e701",
        1412 => x"93d72700",
        1413 => x"b367f800",
        1414 => x"13582740",
        1415 => x"93184800",
        1416 => x"13d3c701",
        1417 => x"33e36800",
        1418 => x"33733301",
        1419 => x"b3f83701",
        1420 => x"135e8801",
        1421 => x"1357f741",
        1422 => x"b3886800",
        1423 => x"b388c801",
        1424 => x"1373d700",
        1425 => x"b3886800",
        1426 => x"b3f84803",
        1427 => x"137727ff",
        1428 => x"939c4700",
        1429 => x"b38cfc40",
        1430 => x"939c2c00",
        1431 => x"b30c9c41",
        1432 => x"b388e800",
        1433 => x"33871741",
        1434 => x"93d8f841",
        1435 => x"33b3e700",
        1436 => x"33081841",
        1437 => x"33086840",
        1438 => x"33082803",
        1439 => x"33035703",
        1440 => x"b3382703",
        1441 => x"33086800",
        1442 => x"33072703",
        1443 => x"33081801",
        1444 => x"9358f841",
        1445 => x"93f83800",
        1446 => x"3387e800",
        1447 => x"b3381701",
        1448 => x"b3880801",
        1449 => x"9398e801",
        1450 => x"13572700",
        1451 => x"33e7e800",
        1452 => x"13184700",
        1453 => x"3307e840",
        1454 => x"13172700",
        1455 => x"338de740",
        1456 => x"eff0cf82",
        1457 => x"83260101",
        1458 => x"13070500",
        1459 => x"13880c00",
        1460 => x"93070d00",
        1461 => x"13060c00",
        1462 => x"93058be5",
        1463 => x"13058101",
        1464 => x"ef00c015",
        1465 => x"13058101",
        1466 => x"efe05ffc",
        1467 => x"e3980be4",
        1468 => x"6ff05fe6",
        1469 => x"03a5c187",
        1470 => x"67800000",
        1471 => x"130101ff",
        1472 => x"23248100",
        1473 => x"23261100",
        1474 => x"93070000",
        1475 => x"13040500",
        1476 => x"63880700",
        1477 => x"93050000",
        1478 => x"97000000",
        1479 => x"e7000000",
        1480 => x"b7370000",
        1481 => x"03a587fb",
        1482 => x"83278502",
        1483 => x"63840700",
        1484 => x"e7800700",
        1485 => x"13050400",
        1486 => x"ef100035",
        1487 => x"130101ff",
        1488 => x"23248100",
        1489 => x"23229100",
        1490 => x"37340000",
        1491 => x"b7340000",
        1492 => x"9387c4fb",
        1493 => x"1304c4fb",
        1494 => x"3304f440",
        1495 => x"23202101",
        1496 => x"23261100",
        1497 => x"13542440",
        1498 => x"9384c4fb",
        1499 => x"13090000",
        1500 => x"63108904",
        1501 => x"b7340000",
        1502 => x"37340000",
        1503 => x"9387c4fb",
        1504 => x"1304c4fb",
        1505 => x"3304f440",
        1506 => x"13542440",
        1507 => x"9384c4fb",
        1508 => x"13090000",
        1509 => x"63188902",
        1510 => x"8320c100",
        1511 => x"03248100",
        1512 => x"83244100",
        1513 => x"03290100",
        1514 => x"13010101",
        1515 => x"67800000",
        1516 => x"83a70400",
        1517 => x"13091900",
        1518 => x"93844400",
        1519 => x"e7800700",
        1520 => x"6ff01ffb",
        1521 => x"83a70400",
        1522 => x"13091900",
        1523 => x"93844400",
        1524 => x"e7800700",
        1525 => x"6ff01ffc",
        1526 => x"130101f6",
        1527 => x"232af108",
        1528 => x"b7070080",
        1529 => x"93c7f7ff",
        1530 => x"232ef100",
        1531 => x"2328f100",
        1532 => x"b707ffff",
        1533 => x"2326d108",
        1534 => x"2324b100",
        1535 => x"232cb100",
        1536 => x"93878720",
        1537 => x"9306c108",
        1538 => x"93058100",
        1539 => x"232e1106",
        1540 => x"232af100",
        1541 => x"2328e108",
        1542 => x"232c0109",
        1543 => x"232e1109",
        1544 => x"2322d100",
        1545 => x"ef00c040",
        1546 => x"83278100",
        1547 => x"23800700",
        1548 => x"8320c107",
        1549 => x"1301010a",
        1550 => x"67800000",
        1551 => x"130101f6",
        1552 => x"232af108",
        1553 => x"b7070080",
        1554 => x"93c7f7ff",
        1555 => x"232ef100",
        1556 => x"2328f100",
        1557 => x"b707ffff",
        1558 => x"93878720",
        1559 => x"232af100",
        1560 => x"2324a100",
        1561 => x"232ca100",
        1562 => x"03a5c187",
        1563 => x"2324c108",
        1564 => x"2326d108",
        1565 => x"13860500",
        1566 => x"93068108",
        1567 => x"93058100",
        1568 => x"232e1106",
        1569 => x"2328e108",
        1570 => x"232c0109",
        1571 => x"232e1109",
        1572 => x"2322d100",
        1573 => x"ef00c039",
        1574 => x"83278100",
        1575 => x"23800700",
        1576 => x"8320c107",
        1577 => x"1301010a",
        1578 => x"67800000",
        1579 => x"13860500",
        1580 => x"93050500",
        1581 => x"03a5c187",
        1582 => x"6f004000",
        1583 => x"130101ff",
        1584 => x"23248100",
        1585 => x"23229100",
        1586 => x"13040500",
        1587 => x"13850500",
        1588 => x"93050600",
        1589 => x"23261100",
        1590 => x"23a20188",
        1591 => x"ef10c01d",
        1592 => x"9307f0ff",
        1593 => x"6318f500",
        1594 => x"83a74188",
        1595 => x"63840700",
        1596 => x"2320f400",
        1597 => x"8320c100",
        1598 => x"03248100",
        1599 => x"83244100",
        1600 => x"13010101",
        1601 => x"67800000",
        1602 => x"130101fe",
        1603 => x"23282101",
        1604 => x"03a98500",
        1605 => x"232c8100",
        1606 => x"23263101",
        1607 => x"23225101",
        1608 => x"23206101",
        1609 => x"232e1100",
        1610 => x"232a9100",
        1611 => x"23244101",
        1612 => x"83aa0500",
        1613 => x"13840500",
        1614 => x"130b0600",
        1615 => x"93890600",
        1616 => x"63ec2609",
        1617 => x"8397c500",
        1618 => x"13f70748",
        1619 => x"63040708",
        1620 => x"03274401",
        1621 => x"93043000",
        1622 => x"83a50501",
        1623 => x"b384e402",
        1624 => x"13072000",
        1625 => x"b38aba40",
        1626 => x"130a0500",
        1627 => x"b3c4e402",
        1628 => x"13871600",
        1629 => x"33075701",
        1630 => x"63f4e400",
        1631 => x"93040700",
        1632 => x"93f70740",
        1633 => x"6386070a",
        1634 => x"93850400",
        1635 => x"13050a00",
        1636 => x"ef001067",
        1637 => x"13090500",
        1638 => x"630c050a",
        1639 => x"83250401",
        1640 => x"13860a00",
        1641 => x"eff05f9d",
        1642 => x"8357c400",
        1643 => x"93f7f7b7",
        1644 => x"93e70708",
        1645 => x"2316f400",
        1646 => x"23282401",
        1647 => x"232a9400",
        1648 => x"33095901",
        1649 => x"b3845441",
        1650 => x"23202401",
        1651 => x"23249400",
        1652 => x"13890900",
        1653 => x"63f42901",
        1654 => x"13890900",
        1655 => x"03250400",
        1656 => x"13060900",
        1657 => x"93050b00",
        1658 => x"eff01f9d",
        1659 => x"83278400",
        1660 => x"13050000",
        1661 => x"b3872741",
        1662 => x"2324f400",
        1663 => x"83270400",
        1664 => x"b3872701",
        1665 => x"2320f400",
        1666 => x"8320c101",
        1667 => x"03248101",
        1668 => x"83244101",
        1669 => x"03290101",
        1670 => x"8329c100",
        1671 => x"032a8100",
        1672 => x"832a4100",
        1673 => x"032b0100",
        1674 => x"13010102",
        1675 => x"67800000",
        1676 => x"13860400",
        1677 => x"13050a00",
        1678 => x"ef001071",
        1679 => x"13090500",
        1680 => x"e31c05f6",
        1681 => x"83250401",
        1682 => x"13050a00",
        1683 => x"ef00d04b",
        1684 => x"9307c000",
        1685 => x"2320fa00",
        1686 => x"8357c400",
        1687 => x"1305f0ff",
        1688 => x"93e70704",
        1689 => x"2316f400",
        1690 => x"6ff01ffa",
        1691 => x"83278600",
        1692 => x"130101fd",
        1693 => x"232e3101",
        1694 => x"23286101",
        1695 => x"23261102",
        1696 => x"23248102",
        1697 => x"23229102",
        1698 => x"23202103",
        1699 => x"232c4101",
        1700 => x"232a5101",
        1701 => x"23267101",
        1702 => x"23248101",
        1703 => x"23229101",
        1704 => x"2320a101",
        1705 => x"032b0600",
        1706 => x"93090600",
        1707 => x"63940712",
        1708 => x"13050000",
        1709 => x"8320c102",
        1710 => x"03248102",
        1711 => x"23a20900",
        1712 => x"83244102",
        1713 => x"03290102",
        1714 => x"8329c101",
        1715 => x"032a8101",
        1716 => x"832a4101",
        1717 => x"032b0101",
        1718 => x"832bc100",
        1719 => x"032c8100",
        1720 => x"832c4100",
        1721 => x"032d0100",
        1722 => x"13010103",
        1723 => x"67800000",
        1724 => x"832b0b00",
        1725 => x"032d4b00",
        1726 => x"130b8b00",
        1727 => x"03298400",
        1728 => x"832a0400",
        1729 => x"e3060dfe",
        1730 => x"63642d09",
        1731 => x"8317c400",
        1732 => x"13f70748",
        1733 => x"630e0706",
        1734 => x"83244401",
        1735 => x"83250401",
        1736 => x"b3049c02",
        1737 => x"b38aba40",
        1738 => x"13871a00",
        1739 => x"3307a701",
        1740 => x"b3c49403",
        1741 => x"63f4e400",
        1742 => x"93040700",
        1743 => x"93f70740",
        1744 => x"6388070a",
        1745 => x"93850400",
        1746 => x"13050a00",
        1747 => x"ef00504b",
        1748 => x"13090500",
        1749 => x"630e050a",
        1750 => x"83250401",
        1751 => x"13860a00",
        1752 => x"eff09f81",
        1753 => x"8357c400",
        1754 => x"93f7f7b7",
        1755 => x"93e70708",
        1756 => x"2316f400",
        1757 => x"23282401",
        1758 => x"232a9400",
        1759 => x"33095901",
        1760 => x"b3845441",
        1761 => x"23202401",
        1762 => x"23249400",
        1763 => x"13090d00",
        1764 => x"63742d01",
        1765 => x"13090d00",
        1766 => x"03250400",
        1767 => x"13060900",
        1768 => x"93850b00",
        1769 => x"eff05f81",
        1770 => x"83278400",
        1771 => x"b3872741",
        1772 => x"2324f400",
        1773 => x"83270400",
        1774 => x"b3872701",
        1775 => x"2320f400",
        1776 => x"83a78900",
        1777 => x"b387a741",
        1778 => x"23a4f900",
        1779 => x"e39207f2",
        1780 => x"6ff01fee",
        1781 => x"130a0500",
        1782 => x"13840500",
        1783 => x"930b0000",
        1784 => x"130d0000",
        1785 => x"130c3000",
        1786 => x"930c2000",
        1787 => x"6ff01ff1",
        1788 => x"13860400",
        1789 => x"13050a00",
        1790 => x"ef001055",
        1791 => x"13090500",
        1792 => x"e31a05f6",
        1793 => x"83250401",
        1794 => x"13050a00",
        1795 => x"ef00d02f",
        1796 => x"9307c000",
        1797 => x"2320fa00",
        1798 => x"8357c400",
        1799 => x"1305f0ff",
        1800 => x"93e70704",
        1801 => x"2316f400",
        1802 => x"23a40900",
        1803 => x"6ff09fe8",
        1804 => x"83d7c500",
        1805 => x"130101f5",
        1806 => x"2324810a",
        1807 => x"2322910a",
        1808 => x"2320210b",
        1809 => x"232c4109",
        1810 => x"2326110a",
        1811 => x"232e3109",
        1812 => x"232a5109",
        1813 => x"23286109",
        1814 => x"23267109",
        1815 => x"23248109",
        1816 => x"23229109",
        1817 => x"2320a109",
        1818 => x"232eb107",
        1819 => x"93f70708",
        1820 => x"130a0500",
        1821 => x"13890500",
        1822 => x"93040600",
        1823 => x"13840600",
        1824 => x"63880706",
        1825 => x"83a70501",
        1826 => x"63940706",
        1827 => x"93050004",
        1828 => x"ef001037",
        1829 => x"2320a900",
        1830 => x"2328a900",
        1831 => x"63160504",
        1832 => x"9307c000",
        1833 => x"2320fa00",
        1834 => x"1305f0ff",
        1835 => x"8320c10a",
        1836 => x"0324810a",
        1837 => x"8324410a",
        1838 => x"0329010a",
        1839 => x"8329c109",
        1840 => x"032a8109",
        1841 => x"832a4109",
        1842 => x"032b0109",
        1843 => x"832bc108",
        1844 => x"032c8108",
        1845 => x"832c4108",
        1846 => x"032d0108",
        1847 => x"832dc107",
        1848 => x"1301010b",
        1849 => x"67800000",
        1850 => x"93070004",
        1851 => x"232af900",
        1852 => x"93070002",
        1853 => x"a304f102",
        1854 => x"93070003",
        1855 => x"23220102",
        1856 => x"2305f102",
        1857 => x"23268100",
        1858 => x"930c5002",
        1859 => x"373b0000",
        1860 => x"b73b0000",
        1861 => x"373d0000",
        1862 => x"372c0000",
        1863 => x"930a0000",
        1864 => x"13840400",
        1865 => x"83470400",
        1866 => x"63840700",
        1867 => x"639c970d",
        1868 => x"b30d9440",
        1869 => x"63069402",
        1870 => x"93860d00",
        1871 => x"13860400",
        1872 => x"93050900",
        1873 => x"13050a00",
        1874 => x"eff01fbc",
        1875 => x"9307f0ff",
        1876 => x"6304f524",
        1877 => x"83274102",
        1878 => x"b387b701",
        1879 => x"2322f102",
        1880 => x"83470400",
        1881 => x"638a0722",
        1882 => x"9307f0ff",
        1883 => x"93041400",
        1884 => x"23280100",
        1885 => x"232e0100",
        1886 => x"232af100",
        1887 => x"232c0100",
        1888 => x"a3090104",
        1889 => x"23240106",
        1890 => x"930d1000",
        1891 => x"83c50400",
        1892 => x"13065000",
        1893 => x"13054bf2",
        1894 => x"ef00d014",
        1895 => x"83270101",
        1896 => x"13841400",
        1897 => x"63140506",
        1898 => x"13f70701",
        1899 => x"63060700",
        1900 => x"13070002",
        1901 => x"a309e104",
        1902 => x"13f78700",
        1903 => x"63060700",
        1904 => x"1307b002",
        1905 => x"a309e104",
        1906 => x"83c60400",
        1907 => x"1307a002",
        1908 => x"638ce604",
        1909 => x"8327c101",
        1910 => x"13840400",
        1911 => x"93060000",
        1912 => x"13069000",
        1913 => x"1305a000",
        1914 => x"03470400",
        1915 => x"93051400",
        1916 => x"130707fd",
        1917 => x"637ee608",
        1918 => x"63840604",
        1919 => x"232ef100",
        1920 => x"6f000004",
        1921 => x"13041400",
        1922 => x"6ff0dff1",
        1923 => x"13074bf2",
        1924 => x"3305e540",
        1925 => x"3395ad00",
        1926 => x"b3e7a700",
        1927 => x"2328f100",
        1928 => x"93040400",
        1929 => x"6ff09ff6",
        1930 => x"0327c100",
        1931 => x"93064700",
        1932 => x"03270700",
        1933 => x"2326d100",
        1934 => x"63420704",
        1935 => x"232ee100",
        1936 => x"03470400",
        1937 => x"9307e002",
        1938 => x"6314f708",
        1939 => x"03471400",
        1940 => x"9307a002",
        1941 => x"6318f704",
        1942 => x"8327c100",
        1943 => x"13042400",
        1944 => x"13874700",
        1945 => x"83a70700",
        1946 => x"2326e100",
        1947 => x"63d40700",
        1948 => x"9307f0ff",
        1949 => x"232af100",
        1950 => x"6f008005",
        1951 => x"3307e040",
        1952 => x"93e72700",
        1953 => x"232ee100",
        1954 => x"2328f100",
        1955 => x"6ff05ffb",
        1956 => x"b387a702",
        1957 => x"13840500",
        1958 => x"93061000",
        1959 => x"b387e700",
        1960 => x"6ff09ff4",
        1961 => x"13041400",
        1962 => x"232a0100",
        1963 => x"93060000",
        1964 => x"93070000",
        1965 => x"13069000",
        1966 => x"1305a000",
        1967 => x"03470400",
        1968 => x"93051400",
        1969 => x"130707fd",
        1970 => x"6372e608",
        1971 => x"e39406fa",
        1972 => x"83450400",
        1973 => x"13063000",
        1974 => x"1385cbf2",
        1975 => x"ef009000",
        1976 => x"63020502",
        1977 => x"9387cbf2",
        1978 => x"3305f540",
        1979 => x"83270101",
        1980 => x"13070004",
        1981 => x"3317a700",
        1982 => x"b3e7e700",
        1983 => x"13041400",
        1984 => x"2328f100",
        1985 => x"83450400",
        1986 => x"13066000",
        1987 => x"13050df3",
        1988 => x"93041400",
        1989 => x"2304b102",
        1990 => x"ef00c07c",
        1991 => x"63080508",
        1992 => x"63980a04",
        1993 => x"03270101",
        1994 => x"8327c100",
        1995 => x"13770710",
        1996 => x"63080702",
        1997 => x"93874700",
        1998 => x"2326f100",
        1999 => x"83274102",
        2000 => x"b3873701",
        2001 => x"2322f102",
        2002 => x"6ff09fdd",
        2003 => x"b387a702",
        2004 => x"13840500",
        2005 => x"93061000",
        2006 => x"b387e700",
        2007 => x"6ff01ff6",
        2008 => x"93877700",
        2009 => x"93f787ff",
        2010 => x"93878700",
        2011 => x"6ff0dffc",
        2012 => x"1307c100",
        2013 => x"93068c90",
        2014 => x"13060900",
        2015 => x"93050101",
        2016 => x"13050a00",
        2017 => x"97000000",
        2018 => x"e7000000",
        2019 => x"9307f0ff",
        2020 => x"93090500",
        2021 => x"e314f5fa",
        2022 => x"8357c900",
        2023 => x"93f70704",
        2024 => x"e39407d0",
        2025 => x"03254102",
        2026 => x"6ff05fd0",
        2027 => x"1307c100",
        2028 => x"93068c90",
        2029 => x"13060900",
        2030 => x"93050101",
        2031 => x"13050a00",
        2032 => x"ef00801b",
        2033 => x"6ff09ffc",
        2034 => x"130101fd",
        2035 => x"232a5101",
        2036 => x"83a70501",
        2037 => x"930a0700",
        2038 => x"03a78500",
        2039 => x"23248102",
        2040 => x"23202103",
        2041 => x"232e3101",
        2042 => x"232c4101",
        2043 => x"23261102",
        2044 => x"23229102",
        2045 => x"23286101",
        2046 => x"23267101",
        2047 => x"93090500",
        2048 => x"13840500",
        2049 => x"13090600",
        2050 => x"138a0600",
        2051 => x"63d4e700",
        2052 => x"93070700",
        2053 => x"2320f900",
        2054 => x"03473404",
        2055 => x"63060700",
        2056 => x"93871700",
        2057 => x"2320f900",
        2058 => x"83270400",
        2059 => x"93f70702",
        2060 => x"63880700",
        2061 => x"83270900",
        2062 => x"93872700",
        2063 => x"2320f900",
        2064 => x"83240400",
        2065 => x"93f46400",
        2066 => x"639e0400",
        2067 => x"130b9401",
        2068 => x"930bf0ff",
        2069 => x"8327c400",
        2070 => x"03270900",
        2071 => x"b387e740",
        2072 => x"63c2f408",
        2073 => x"83473404",
        2074 => x"b336f000",
        2075 => x"83270400",
        2076 => x"93f70702",
        2077 => x"6390070c",
        2078 => x"13063404",
        2079 => x"93050a00",
        2080 => x"13850900",
        2081 => x"e7800a00",
        2082 => x"9307f0ff",
        2083 => x"6308f506",
        2084 => x"83270400",
        2085 => x"13074000",
        2086 => x"93040000",
        2087 => x"93f76700",
        2088 => x"639ce700",
        2089 => x"8324c400",
        2090 => x"83270900",
        2091 => x"b384f440",
        2092 => x"63d40400",
        2093 => x"93040000",
        2094 => x"83278400",
        2095 => x"03270401",
        2096 => x"6356f700",
        2097 => x"b387e740",
        2098 => x"b384f400",
        2099 => x"13090000",
        2100 => x"1304a401",
        2101 => x"130bf0ff",
        2102 => x"63902409",
        2103 => x"13050000",
        2104 => x"6f000002",
        2105 => x"93061000",
        2106 => x"13060b00",
        2107 => x"93050a00",
        2108 => x"13850900",
        2109 => x"e7800a00",
        2110 => x"631a7503",
        2111 => x"1305f0ff",
        2112 => x"8320c102",
        2113 => x"03248102",
        2114 => x"83244102",
        2115 => x"03290102",
        2116 => x"8329c101",
        2117 => x"032a8101",
        2118 => x"832a4101",
        2119 => x"032b0101",
        2120 => x"832bc100",
        2121 => x"13010103",
        2122 => x"67800000",
        2123 => x"93841400",
        2124 => x"6ff05ff2",
        2125 => x"3307d400",
        2126 => x"13060003",
        2127 => x"a301c704",
        2128 => x"03475404",
        2129 => x"93871600",
        2130 => x"b307f400",
        2131 => x"93862600",
        2132 => x"a381e704",
        2133 => x"6ff05ff2",
        2134 => x"93061000",
        2135 => x"13060400",
        2136 => x"93050a00",
        2137 => x"13850900",
        2138 => x"e7800a00",
        2139 => x"e30865f9",
        2140 => x"13091900",
        2141 => x"6ff05ff6",
        2142 => x"130101fd",
        2143 => x"23248102",
        2144 => x"23229102",
        2145 => x"23202103",
        2146 => x"232e3101",
        2147 => x"23261102",
        2148 => x"232c4101",
        2149 => x"232a5101",
        2150 => x"23286101",
        2151 => x"83c88501",
        2152 => x"93078007",
        2153 => x"93040500",
        2154 => x"13840500",
        2155 => x"13090600",
        2156 => x"93890600",
        2157 => x"63ee1701",
        2158 => x"93072006",
        2159 => x"93863504",
        2160 => x"63ee1701",
        2161 => x"638a082a",
        2162 => x"93078005",
        2163 => x"638af820",
        2164 => x"930a2404",
        2165 => x"23011405",
        2166 => x"6f004004",
        2167 => x"9387d8f9",
        2168 => x"93f7f70f",
        2169 => x"13065001",
        2170 => x"e364f6fe",
        2171 => x"37360000",
        2172 => x"93972700",
        2173 => x"130606f6",
        2174 => x"b387c700",
        2175 => x"83a70700",
        2176 => x"67800700",
        2177 => x"83270700",
        2178 => x"938a2504",
        2179 => x"93864700",
        2180 => x"83a70700",
        2181 => x"2320d700",
        2182 => x"2381f504",
        2183 => x"93071000",
        2184 => x"6f004029",
        2185 => x"03a60500",
        2186 => x"83270700",
        2187 => x"13750608",
        2188 => x"93854700",
        2189 => x"630e0504",
        2190 => x"83a70700",
        2191 => x"2320b700",
        2192 => x"37370000",
        2193 => x"83254400",
        2194 => x"130887f3",
        2195 => x"63d2071e",
        2196 => x"1307d002",
        2197 => x"a301e404",
        2198 => x"2324b400",
        2199 => x"63d80504",
        2200 => x"b307f040",
        2201 => x"1307a000",
        2202 => x"938a0600",
        2203 => x"33f6e702",
        2204 => x"938afaff",
        2205 => x"3306c800",
        2206 => x"03460600",
        2207 => x"2380ca00",
        2208 => x"13860700",
        2209 => x"b3d7e702",
        2210 => x"e372e6fe",
        2211 => x"6f008009",
        2212 => x"83a70700",
        2213 => x"13750604",
        2214 => x"2320b700",
        2215 => x"e30205fa",
        2216 => x"93970701",
        2217 => x"93d70741",
        2218 => x"6ff09ff9",
        2219 => x"1376b6ff",
        2220 => x"2320c400",
        2221 => x"6ff0dffa",
        2222 => x"03a60500",
        2223 => x"83270700",
        2224 => x"13750608",
        2225 => x"93854700",
        2226 => x"63080500",
        2227 => x"2320b700",
        2228 => x"83a70700",
        2229 => x"6f004001",
        2230 => x"13760604",
        2231 => x"2320b700",
        2232 => x"e30806fe",
        2233 => x"83d70700",
        2234 => x"37380000",
        2235 => x"1307f006",
        2236 => x"130888f3",
        2237 => x"639ae812",
        2238 => x"13078000",
        2239 => x"a3010404",
        2240 => x"03264400",
        2241 => x"2324c400",
        2242 => x"e34006f6",
        2243 => x"83250400",
        2244 => x"93f5b5ff",
        2245 => x"2320b400",
        2246 => x"e39807f4",
        2247 => x"938a0600",
        2248 => x"e31406f4",
        2249 => x"93078000",
        2250 => x"6314f702",
        2251 => x"83270400",
        2252 => x"93f71700",
        2253 => x"638e0700",
        2254 => x"03274400",
        2255 => x"83270401",
        2256 => x"63c8e700",
        2257 => x"93070003",
        2258 => x"a38ffafe",
        2259 => x"938afaff",
        2260 => x"b3865641",
        2261 => x"2328d400",
        2262 => x"13870900",
        2263 => x"93060900",
        2264 => x"1306c100",
        2265 => x"93050400",
        2266 => x"13850400",
        2267 => x"eff0dfc5",
        2268 => x"130af0ff",
        2269 => x"63164515",
        2270 => x"1305f0ff",
        2271 => x"8320c102",
        2272 => x"03248102",
        2273 => x"83244102",
        2274 => x"03290102",
        2275 => x"8329c101",
        2276 => x"032a8101",
        2277 => x"832a4101",
        2278 => x"032b0101",
        2279 => x"13010103",
        2280 => x"67800000",
        2281 => x"83a70500",
        2282 => x"93e70702",
        2283 => x"23a0f500",
        2284 => x"37380000",
        2285 => x"93088007",
        2286 => x"1308c8f4",
        2287 => x"03260400",
        2288 => x"a3021405",
        2289 => x"83270700",
        2290 => x"13750608",
        2291 => x"93854700",
        2292 => x"630e0500",
        2293 => x"2320b700",
        2294 => x"83a70700",
        2295 => x"6f000002",
        2296 => x"37380000",
        2297 => x"130888f3",
        2298 => x"6ff05ffd",
        2299 => x"13750604",
        2300 => x"2320b700",
        2301 => x"e30205fe",
        2302 => x"83d70700",
        2303 => x"13771600",
        2304 => x"63060700",
        2305 => x"13660602",
        2306 => x"2320c400",
        2307 => x"63860700",
        2308 => x"13070001",
        2309 => x"6ff09fee",
        2310 => x"03270400",
        2311 => x"1377f7fd",
        2312 => x"2320e400",
        2313 => x"6ff0dffe",
        2314 => x"1307a000",
        2315 => x"6ff01fed",
        2316 => x"130887f3",
        2317 => x"1307a000",
        2318 => x"6ff09fec",
        2319 => x"03a60500",
        2320 => x"83270700",
        2321 => x"83a54501",
        2322 => x"13780608",
        2323 => x"13854700",
        2324 => x"630a0800",
        2325 => x"2320a700",
        2326 => x"83a70700",
        2327 => x"23a0b700",
        2328 => x"6f008001",
        2329 => x"2320a700",
        2330 => x"13760604",
        2331 => x"83a70700",
        2332 => x"e30606fe",
        2333 => x"2390b700",
        2334 => x"23280400",
        2335 => x"938a0600",
        2336 => x"6ff09fed",
        2337 => x"83270700",
        2338 => x"03a64500",
        2339 => x"93050000",
        2340 => x"93864700",
        2341 => x"2320d700",
        2342 => x"83aa0700",
        2343 => x"13850a00",
        2344 => x"ef004024",
        2345 => x"63060500",
        2346 => x"33055541",
        2347 => x"2322a400",
        2348 => x"83274400",
        2349 => x"2328f400",
        2350 => x"a3010404",
        2351 => x"6ff0dfe9",
        2352 => x"83260401",
        2353 => x"13860a00",
        2354 => x"93050900",
        2355 => x"13850400",
        2356 => x"e7800900",
        2357 => x"e30245eb",
        2358 => x"83270400",
        2359 => x"93f72700",
        2360 => x"63940704",
        2361 => x"8327c100",
        2362 => x"0325c400",
        2363 => x"e358f5e8",
        2364 => x"13850700",
        2365 => x"6ff09fe8",
        2366 => x"93061000",
        2367 => x"13860a00",
        2368 => x"93050900",
        2369 => x"13850400",
        2370 => x"e7800900",
        2371 => x"e30665e7",
        2372 => x"130a1a00",
        2373 => x"8327c400",
        2374 => x"0327c100",
        2375 => x"b387e740",
        2376 => x"e34cfafc",
        2377 => x"6ff01ffc",
        2378 => x"130a0000",
        2379 => x"930a9401",
        2380 => x"130bf0ff",
        2381 => x"6ff01ffe",
        2382 => x"130101ff",
        2383 => x"23248100",
        2384 => x"13840500",
        2385 => x"83a50500",
        2386 => x"23229100",
        2387 => x"23261100",
        2388 => x"93040500",
        2389 => x"63840500",
        2390 => x"eff01ffe",
        2391 => x"93050400",
        2392 => x"03248100",
        2393 => x"8320c100",
        2394 => x"13850400",
        2395 => x"83244100",
        2396 => x"13010101",
        2397 => x"6f004019",
        2398 => x"83a7c187",
        2399 => x"6382a716",
        2400 => x"83274502",
        2401 => x"130101fe",
        2402 => x"232c8100",
        2403 => x"232e1100",
        2404 => x"232a9100",
        2405 => x"23282101",
        2406 => x"23263101",
        2407 => x"13040500",
        2408 => x"638a0704",
        2409 => x"83a7c700",
        2410 => x"638c0702",
        2411 => x"93040000",
        2412 => x"13090008",
        2413 => x"83274402",
        2414 => x"83a7c700",
        2415 => x"b3879700",
        2416 => x"83a50700",
        2417 => x"6396050e",
        2418 => x"93844400",
        2419 => x"e39424ff",
        2420 => x"83274402",
        2421 => x"13050400",
        2422 => x"83a5c700",
        2423 => x"ef00c012",
        2424 => x"83274402",
        2425 => x"83a50700",
        2426 => x"63860500",
        2427 => x"13050400",
        2428 => x"ef008011",
        2429 => x"83254401",
        2430 => x"63860500",
        2431 => x"13050400",
        2432 => x"ef008010",
        2433 => x"83254402",
        2434 => x"63860500",
        2435 => x"13050400",
        2436 => x"ef00800f",
        2437 => x"83258403",
        2438 => x"63860500",
        2439 => x"13050400",
        2440 => x"ef00800e",
        2441 => x"8325c403",
        2442 => x"63860500",
        2443 => x"13050400",
        2444 => x"ef00800d",
        2445 => x"83250404",
        2446 => x"63860500",
        2447 => x"13050400",
        2448 => x"ef00800c",
        2449 => x"8325c405",
        2450 => x"63860500",
        2451 => x"13050400",
        2452 => x"ef00800b",
        2453 => x"83258405",
        2454 => x"63860500",
        2455 => x"13050400",
        2456 => x"ef00800a",
        2457 => x"83254403",
        2458 => x"63860500",
        2459 => x"13050400",
        2460 => x"ef008009",
        2461 => x"83278401",
        2462 => x"63860704",
        2463 => x"83278402",
        2464 => x"13050400",
        2465 => x"e7800700",
        2466 => x"83258404",
        2467 => x"638c0502",
        2468 => x"13050400",
        2469 => x"03248101",
        2470 => x"8320c101",
        2471 => x"83244101",
        2472 => x"03290101",
        2473 => x"8329c100",
        2474 => x"13010102",
        2475 => x"6ff0dfe8",
        2476 => x"83a90500",
        2477 => x"13050400",
        2478 => x"ef000005",
        2479 => x"93850900",
        2480 => x"6ff05ff0",
        2481 => x"8320c101",
        2482 => x"03248101",
        2483 => x"83244101",
        2484 => x"03290101",
        2485 => x"8329c100",
        2486 => x"13010102",
        2487 => x"67800000",
        2488 => x"67800000",
        2489 => x"93f5f50f",
        2490 => x"3306c500",
        2491 => x"6316c500",
        2492 => x"13050000",
        2493 => x"67800000",
        2494 => x"83470500",
        2495 => x"e38cb7fe",
        2496 => x"13051500",
        2497 => x"6ff09ffe",
        2498 => x"638a050e",
        2499 => x"83a7c5ff",
        2500 => x"130101fe",
        2501 => x"232c8100",
        2502 => x"232e1100",
        2503 => x"1384c5ff",
        2504 => x"63d40700",
        2505 => x"3304f400",
        2506 => x"2326a100",
        2507 => x"ef008033",
        2508 => x"83a7c188",
        2509 => x"0325c100",
        2510 => x"639e0700",
        2511 => x"23220400",
        2512 => x"23a68188",
        2513 => x"03248101",
        2514 => x"8320c101",
        2515 => x"13010102",
        2516 => x"6f008031",
        2517 => x"6374f402",
        2518 => x"03260400",
        2519 => x"b306c400",
        2520 => x"639ad700",
        2521 => x"83a60700",
        2522 => x"83a74700",
        2523 => x"b386c600",
        2524 => x"2320d400",
        2525 => x"2322f400",
        2526 => x"6ff09ffc",
        2527 => x"13870700",
        2528 => x"83a74700",
        2529 => x"63840700",
        2530 => x"e37af4fe",
        2531 => x"83260700",
        2532 => x"3306d700",
        2533 => x"63188602",
        2534 => x"03260400",
        2535 => x"b386c600",
        2536 => x"2320d700",
        2537 => x"3306d700",
        2538 => x"e39ec7f8",
        2539 => x"03a60700",
        2540 => x"83a74700",
        2541 => x"b306d600",
        2542 => x"2320d700",
        2543 => x"2322f700",
        2544 => x"6ff05ff8",
        2545 => x"6378c400",
        2546 => x"9307c000",
        2547 => x"2320f500",
        2548 => x"6ff05ff7",
        2549 => x"03260400",
        2550 => x"b306c400",
        2551 => x"639ad700",
        2552 => x"83a60700",
        2553 => x"83a74700",
        2554 => x"b386c600",
        2555 => x"2320d400",
        2556 => x"2322f400",
        2557 => x"23228700",
        2558 => x"6ff0dff4",
        2559 => x"67800000",
        2560 => x"130101fe",
        2561 => x"232a9100",
        2562 => x"93843500",
        2563 => x"93f4c4ff",
        2564 => x"23282101",
        2565 => x"232e1100",
        2566 => x"232c8100",
        2567 => x"23263101",
        2568 => x"93848400",
        2569 => x"9307c000",
        2570 => x"13090500",
        2571 => x"63f0f406",
        2572 => x"9304c000",
        2573 => x"63eeb404",
        2574 => x"13050900",
        2575 => x"ef008022",
        2576 => x"03a7c188",
        2577 => x"13040700",
        2578 => x"63180406",
        2579 => x"83a78188",
        2580 => x"639a0700",
        2581 => x"93050000",
        2582 => x"13050900",
        2583 => x"ef00001c",
        2584 => x"23a4a188",
        2585 => x"93850400",
        2586 => x"13050900",
        2587 => x"ef00001b",
        2588 => x"9309f0ff",
        2589 => x"631a350b",
        2590 => x"9307c000",
        2591 => x"2320f900",
        2592 => x"13050900",
        2593 => x"ef00401e",
        2594 => x"6f000001",
        2595 => x"e3d404fa",
        2596 => x"9307c000",
        2597 => x"2320f900",
        2598 => x"13050000",
        2599 => x"8320c101",
        2600 => x"03248101",
        2601 => x"83244101",
        2602 => x"03290101",
        2603 => x"8329c100",
        2604 => x"13010102",
        2605 => x"67800000",
        2606 => x"83270400",
        2607 => x"b3879740",
        2608 => x"63ce0704",
        2609 => x"1306b000",
        2610 => x"637af600",
        2611 => x"2320f400",
        2612 => x"3304f400",
        2613 => x"23209400",
        2614 => x"6f000001",
        2615 => x"83274400",
        2616 => x"631a8702",
        2617 => x"23a6f188",
        2618 => x"13050900",
        2619 => x"ef00c017",
        2620 => x"1305b400",
        2621 => x"93074400",
        2622 => x"137585ff",
        2623 => x"3307f540",
        2624 => x"e30ef5f8",
        2625 => x"3304e400",
        2626 => x"b387a740",
        2627 => x"2320f400",
        2628 => x"6ff0dff8",
        2629 => x"2322f700",
        2630 => x"6ff01ffd",
        2631 => x"13070400",
        2632 => x"03244400",
        2633 => x"6ff05ff2",
        2634 => x"13043500",
        2635 => x"1374c4ff",
        2636 => x"e30285fa",
        2637 => x"b305a440",
        2638 => x"13050900",
        2639 => x"ef00000e",
        2640 => x"e31a35f9",
        2641 => x"6ff05ff3",
        2642 => x"130101fe",
        2643 => x"232c8100",
        2644 => x"232e1100",
        2645 => x"232a9100",
        2646 => x"23282101",
        2647 => x"23263101",
        2648 => x"23244101",
        2649 => x"13040600",
        2650 => x"63940502",
        2651 => x"03248101",
        2652 => x"8320c101",
        2653 => x"83244101",
        2654 => x"03290101",
        2655 => x"8329c100",
        2656 => x"032a8100",
        2657 => x"93050600",
        2658 => x"13010102",
        2659 => x"6ff05fe7",
        2660 => x"63180602",
        2661 => x"eff05fd7",
        2662 => x"93040000",
        2663 => x"8320c101",
        2664 => x"03248101",
        2665 => x"03290101",
        2666 => x"8329c100",
        2667 => x"032a8100",
        2668 => x"13850400",
        2669 => x"83244101",
        2670 => x"13010102",
        2671 => x"67800000",
        2672 => x"130a0500",
        2673 => x"93840500",
        2674 => x"ef00400a",
        2675 => x"13090500",
        2676 => x"63668500",
        2677 => x"93571500",
        2678 => x"e3e287fc",
        2679 => x"93050400",
        2680 => x"13050a00",
        2681 => x"eff0dfe1",
        2682 => x"93090500",
        2683 => x"e30605fa",
        2684 => x"13060400",
        2685 => x"63748900",
        2686 => x"13060900",
        2687 => x"93850400",
        2688 => x"13850900",
        2689 => x"efe05f97",
        2690 => x"93850400",
        2691 => x"13050a00",
        2692 => x"eff09fcf",
        2693 => x"93840900",
        2694 => x"6ff05ff8",
        2695 => x"130101ff",
        2696 => x"23248100",
        2697 => x"23229100",
        2698 => x"13040500",
        2699 => x"13850500",
        2700 => x"23261100",
        2701 => x"23a20188",
        2702 => x"ef00000c",
        2703 => x"9307f0ff",
        2704 => x"6318f500",
        2705 => x"83a74188",
        2706 => x"63840700",
        2707 => x"2320f400",
        2708 => x"8320c100",
        2709 => x"03248100",
        2710 => x"83244100",
        2711 => x"13010101",
        2712 => x"67800000",
        2713 => x"67800000",
        2714 => x"67800000",
        2715 => x"83a7c5ff",
        2716 => x"1385c7ff",
        2717 => x"63d80700",
        2718 => x"b385a500",
        2719 => x"83a70500",
        2720 => x"3305f500",
        2721 => x"67800000",
        2722 => x"9308d005",
        2723 => x"73000000",
        2724 => x"63520502",
        2725 => x"130101ff",
        2726 => x"23248100",
        2727 => x"13040500",
        2728 => x"23261100",
        2729 => x"33048040",
        2730 => x"efe0dfc4",
        2731 => x"23208500",
        2732 => x"6f000000",
        2733 => x"6f000000",
        2734 => x"130101ff",
        2735 => x"23261100",
        2736 => x"23248100",
        2737 => x"9308900a",
        2738 => x"73000000",
        2739 => x"13040500",
        2740 => x"635a0500",
        2741 => x"33048040",
        2742 => x"efe0dfc1",
        2743 => x"23208500",
        2744 => x"1304f0ff",
        2745 => x"8320c100",
        2746 => x"13050400",
        2747 => x"03248100",
        2748 => x"13010101",
        2749 => x"67800000",
        2750 => x"03a70189",
        2751 => x"130101ff",
        2752 => x"23261100",
        2753 => x"93070500",
        2754 => x"631c0702",
        2755 => x"9308600d",
        2756 => x"13050000",
        2757 => x"73000000",
        2758 => x"1307f0ff",
        2759 => x"6310e502",
        2760 => x"efe05fbd",
        2761 => x"9307c000",
        2762 => x"2320f500",
        2763 => x"1305f0ff",
        2764 => x"8320c100",
        2765 => x"13010101",
        2766 => x"67800000",
        2767 => x"23a8a188",
        2768 => x"03a70189",
        2769 => x"9308600d",
        2770 => x"b387e700",
        2771 => x"13850700",
        2772 => x"73000000",
        2773 => x"e316f5fc",
        2774 => x"23a8a188",
        2775 => x"13050700",
        2776 => x"6ff01ffd",
        2777 => x"10000000",
        2778 => x"00000000",
        2779 => x"037a5200",
        2780 => x"017c0101",
        2781 => x"1b0d0200",
        2782 => x"10000000",
        2783 => x"18000000",
        2784 => x"6cdbffff",
        2785 => x"78040000",
        2786 => x"00000000",
        2787 => x"10000000",
        2788 => x"00000000",
        2789 => x"037a5200",
        2790 => x"017c0101",
        2791 => x"1b0d0200",
        2792 => x"10000000",
        2793 => x"18000000",
        2794 => x"bcdfffff",
        2795 => x"30040000",
        2796 => x"00000000",
        2797 => x"10000000",
        2798 => x"00000000",
        2799 => x"037a5200",
        2800 => x"017c0101",
        2801 => x"1b0d0200",
        2802 => x"10000000",
        2803 => x"18000000",
        2804 => x"c4e3ffff",
        2805 => x"e4030000",
        2806 => x"00000000",
        2807 => x"30313233",
        2808 => x"34353637",
        2809 => x"38396162",
        2810 => x"63646566",
        2811 => x"00000000",
        2812 => x"44040000",
        2813 => x"50040000",
        2814 => x"20040000",
        2815 => x"38040000",
        2816 => x"2c040000",
        2817 => x"74030000",
        2818 => x"74030000",
        2819 => x"74030000",
        2820 => x"94040000",
        2821 => x"74030000",
        2822 => x"74030000",
        2823 => x"74030000",
        2824 => x"74030000",
        2825 => x"74030000",
        2826 => x"74030000",
        2827 => x"74030000",
        2828 => x"5c040000",
        2829 => x"f8040000",
        2830 => x"b0040000",
        2831 => x"b0040000",
        2832 => x"b0040000",
        2833 => x"b0040000",
        2834 => x"ec040000",
        2835 => x"38050000",
        2836 => x"10050000",
        2837 => x"b0040000",
        2838 => x"b0040000",
        2839 => x"b0040000",
        2840 => x"b0040000",
        2841 => x"b0040000",
        2842 => x"b0040000",
        2843 => x"b0040000",
        2844 => x"b0040000",
        2845 => x"b0040000",
        2846 => x"b0040000",
        2847 => x"b0040000",
        2848 => x"b0040000",
        2849 => x"b0040000",
        2850 => x"b0040000",
        2851 => x"d8040000",
        2852 => x"d8040000",
        2853 => x"b0040000",
        2854 => x"b0040000",
        2855 => x"b0040000",
        2856 => x"b0040000",
        2857 => x"b0040000",
        2858 => x"b0040000",
        2859 => x"b0040000",
        2860 => x"b0040000",
        2861 => x"b0040000",
        2862 => x"b0040000",
        2863 => x"b0040000",
        2864 => x"b0040000",
        2865 => x"ec040000",
        2866 => x"f8040000",
        2867 => x"b4050000",
        2868 => x"9c050000",
        2869 => x"b0040000",
        2870 => x"b0040000",
        2871 => x"b0040000",
        2872 => x"b0040000",
        2873 => x"b0040000",
        2874 => x"b0040000",
        2875 => x"84050000",
        2876 => x"b0040000",
        2877 => x"b0040000",
        2878 => x"b0040000",
        2879 => x"b0040000",
        2880 => x"d8040000",
        2881 => x"d8040000",
        2882 => x"00010202",
        2883 => x"03030303",
        2884 => x"04040404",
        2885 => x"04040404",
        2886 => x"05050505",
        2887 => x"05050505",
        2888 => x"05050505",
        2889 => x"05050505",
        2890 => x"06060606",
        2891 => x"06060606",
        2892 => x"06060606",
        2893 => x"06060606",
        2894 => x"06060606",
        2895 => x"06060606",
        2896 => x"06060606",
        2897 => x"06060606",
        2898 => x"07070707",
        2899 => x"07070707",
        2900 => x"07070707",
        2901 => x"07070707",
        2902 => x"07070707",
        2903 => x"07070707",
        2904 => x"07070707",
        2905 => x"07070707",
        2906 => x"07070707",
        2907 => x"07070707",
        2908 => x"07070707",
        2909 => x"07070707",
        2910 => x"07070707",
        2911 => x"07070707",
        2912 => x"07070707",
        2913 => x"07070707",
        2914 => x"08080808",
        2915 => x"08080808",
        2916 => x"08080808",
        2917 => x"08080808",
        2918 => x"08080808",
        2919 => x"08080808",
        2920 => x"08080808",
        2921 => x"08080808",
        2922 => x"08080808",
        2923 => x"08080808",
        2924 => x"08080808",
        2925 => x"08080808",
        2926 => x"08080808",
        2927 => x"08080808",
        2928 => x"08080808",
        2929 => x"08080808",
        2930 => x"08080808",
        2931 => x"08080808",
        2932 => x"08080808",
        2933 => x"08080808",
        2934 => x"08080808",
        2935 => x"08080808",
        2936 => x"08080808",
        2937 => x"08080808",
        2938 => x"08080808",
        2939 => x"08080808",
        2940 => x"08080808",
        2941 => x"08080808",
        2942 => x"08080808",
        2943 => x"08080808",
        2944 => x"08080808",
        2945 => x"08080808",
        2946 => x"0d0a4542",
        2947 => x"5245414b",
        2948 => x"21206d65",
        2949 => x"7063203d",
        2950 => x"20000000",
        2951 => x"20696e73",
        2952 => x"6e203d20",
        2953 => x"00000000",
        2954 => x"0d0a0d0a",
        2955 => x"44697370",
        2956 => x"6c617969",
        2957 => x"6e672074",
        2958 => x"68652074",
        2959 => x"696d6520",
        2960 => x"70617373",
        2961 => x"65642073",
        2962 => x"696e6365",
        2963 => x"20726573",
        2964 => x"65740d0a",
        2965 => x"0d0a0000",
        2966 => x"2530356c",
        2967 => x"643a2530",
        2968 => x"366c6420",
        2969 => x"20202530",
        2970 => x"326c643a",
        2971 => x"2530326c",
        2972 => x"643a2530",
        2973 => x"326c640d",
        2974 => x"00000000",
        2975 => x"696e7465",
        2976 => x"72727570",
        2977 => x"745f6469",
        2978 => x"72656374",
        2979 => x"00000000",
        2980 => x"54485541",
        2981 => x"53205249",
        2982 => x"53432d56",
        2983 => x"20525633",
        2984 => x"32494d20",
        2985 => x"62617265",
        2986 => x"206d6574",
        2987 => x"616c2070",
        2988 => x"726f6365",
        2989 => x"73736f72",
        2990 => x"00000000",
        2991 => x"54686520",
        2992 => x"48616775",
        2993 => x"6520556e",
        2994 => x"69766572",
        2995 => x"73697479",
        2996 => x"206f6620",
        2997 => x"4170706c",
        2998 => x"69656420",
        2999 => x"53636965",
        3000 => x"6e636573",
        3001 => x"00000000",
        3002 => x"44657061",
        3003 => x"72746d65",
        3004 => x"6e74206f",
        3005 => x"6620456c",
        3006 => x"65637472",
        3007 => x"6963616c",
        3008 => x"20456e67",
        3009 => x"696e6565",
        3010 => x"72696e67",
        3011 => x"00000000",
        3012 => x"4a2e452e",
        3013 => x"4a2e206f",
        3014 => x"70206465",
        3015 => x"6e204272",
        3016 => x"6f757700",
        3017 => x"232d302b",
        3018 => x"20000000",
        3019 => x"686c4c00",
        3020 => x"65666745",
        3021 => x"46470000",
        3022 => x"30313233",
        3023 => x"34353637",
        3024 => x"38394142",
        3025 => x"43444546",
        3026 => x"00000000",
        3027 => x"30313233",
        3028 => x"34353637",
        3029 => x"38396162",
        3030 => x"63646566",
        3031 => x"00000000",
        3032 => x"04220000",
        3033 => x"24220000",
        3034 => x"d0210000",
        3035 => x"d0210000",
        3036 => x"d0210000",
        3037 => x"d0210000",
        3038 => x"24220000",
        3039 => x"d0210000",
        3040 => x"d0210000",
        3041 => x"d0210000",
        3042 => x"d0210000",
        3043 => x"3c240000",
        3044 => x"b8220000",
        3045 => x"a4230000",
        3046 => x"d0210000",
        3047 => x"d0210000",
        3048 => x"84240000",
        3049 => x"d0210000",
        3050 => x"b8220000",
        3051 => x"d0210000",
        3052 => x"d0210000",
        3053 => x"b0230000",
        3054 => x"18000020",
        3055 => x"7c2e0000",
        3056 => x"902e0000",
        3057 => x"bc2e0000",
        3058 => x"e82e0000",
        3059 => x"102f0000",
        3060 => x"00000000",
        3061 => x"00000000",
        3062 => x"00000000",
        3063 => x"00000000",
        3064 => x"00000000",
        3065 => x"00000000",
        3066 => x"00000000",
        3067 => x"00000000",
        3068 => x"00000000",
        3069 => x"00000000",
        3070 => x"00000000",
        3071 => x"00000000",
        3072 => x"00000000",
        3073 => x"00000000",
        3074 => x"00000000",
        3075 => x"00000000",
        3076 => x"00000000",
        3077 => x"00000000",
        3078 => x"00000000",
        3079 => x"00000000",
        3080 => x"00000000",
        3081 => x"00000000",
        3082 => x"00000000",
        3083 => x"00000000",
        3084 => x"00000000",
        3085 => x"80000020",
        3086 => x"18000020",
        others => (others => '0')
    );
end package processor_common_rom;
