-- #################################################################################################
-- # bootloader.vhd - The bootloader ROM                                                           #
-- # ********************************************************************************************* #
-- # This file is part of the THUAS RISCV RV32 Project                                             #
-- # ********************************************************************************************* #
-- # BSD 3-Clause License                                                                          #
-- #                                                                                               #
-- # Copyright (c) 2023, Jesse op den Brouw. All rights reserved.                                  #
-- #                                                                                               #
-- # Redistribution and use in source and binary forms, with or without modification, are          #
-- # permitted provided that the following conditions are met:                                     #
-- #                                                                                               #
-- # 1. Redistributions of source code must retain the above copyright notice, this list of        #
-- #    conditions and the following disclaimer.                                                   #
-- #                                                                                               #
-- # 2. Redistributions in binary form must reproduce the above copyright notice, this list of     #
-- #    conditions and the following disclaimer in the documentation and/or other materials        #
-- #    provided with the distribution.                                                            #
-- #                                                                                               #
-- # 3. Neither the name of the copyright holder nor the names of its contributors may be used to  #
-- #    endorse or promote products derived from this software without specific prior written      #
-- #    permission.                                                                                #
-- #                                                                                               #
-- # THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND ANY EXPRESS   #
-- # OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED WARRANTIES OF               #
-- # MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE    #
-- # COPYRIGHT HOLDER OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL,     #
-- # EXEMPLARY, OR CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE #
-- # GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER CAUSED    #
-- # AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT (INCLUDING     #
-- # NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED  #
-- # OF THE POSSIBILITY OF SUCH DAMAGE.                                                            #
-- # ********************************************************************************************* #
-- # https:/github.com/jesseopdenbrouw/riscv-rv32                                                  #
-- #################################################################################################

-- This file contains the description of the bootloader ROM. The ROM
-- is placed in immutable onboard RAM blocks. A read takes two
-- clock cycles, for both instruction and data.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.processor_common.all;
use work.processor_common_rom.all;

entity bootloader is
    port (I_clk : in std_logic;
          I_areset : in std_logic;
          I_pc : in data_type;
          I_memaddress : in data_type;
          I_memsize : in memsize_type;
          I_csboot : in std_logic;
          I_stall : in std_logic;
          O_instr : out data_type;
          O_dataout : out data_type;
          --
          O_load_misaligned_error : out std_logic
         );
end entity bootloader;

architecture rtl of bootloader is

-- The bootloader ROM
signal bootrom : bootloader_type := (
           0 => x"97020000",
           1 => x"93820208",
           2 => x"73905230",
           3 => x"97010010",
           4 => x"9381417f",
           5 => x"17810010",
           6 => x"1301c1fe",
           7 => x"9387c187",
           8 => x"1387c187",
           9 => x"13060000",
          10 => x"63e4e700",
          11 => x"3386e740",
          12 => x"93050000",
          13 => x"1385c187",
          14 => x"ef000007",
          15 => x"37050020",
          16 => x"9387c187",
          17 => x"13070500",
          18 => x"13060000",
          19 => x"63e4e700",
          20 => x"3386e740",
          21 => x"b7150010",
          22 => x"9385c5f1",
          23 => x"13050500",
          24 => x"ef004002",
          25 => x"ef001026",
          26 => x"b7050020",
          27 => x"13060000",
          28 => x"93850500",
          29 => x"13055000",
          30 => x"ef00c051",
          31 => x"ef009020",
          32 => x"6f000000",
          33 => x"13030500",
          34 => x"630e0600",
          35 => x"83830500",
          36 => x"23007300",
          37 => x"1306f6ff",
          38 => x"13031300",
          39 => x"93851500",
          40 => x"e31606fe",
          41 => x"67800000",
          42 => x"13030500",
          43 => x"630a0600",
          44 => x"2300b300",
          45 => x"1306f6ff",
          46 => x"13031300",
          47 => x"e31a06fe",
          48 => x"67800000",
          49 => x"03460500",
          50 => x"83c60500",
          51 => x"13051500",
          52 => x"93851500",
          53 => x"6314d600",
          54 => x"e31606fe",
          55 => x"3305d640",
          56 => x"67800000",
          57 => x"6f000000",
          58 => x"b70700f0",
          59 => x"03a54702",
          60 => x"13754500",
          61 => x"67800000",
          62 => x"370700f0",
          63 => x"83274702",
          64 => x"93f74700",
          65 => x"e38c07fe",
          66 => x"03258702",
          67 => x"1375f50f",
          68 => x"67800000",
          69 => x"130101fd",
          70 => x"23202103",
          71 => x"37190010",
          72 => x"23248102",
          73 => x"23229102",
          74 => x"232e3101",
          75 => x"232c4101",
          76 => x"232a5101",
          77 => x"23286101",
          78 => x"23267101",
          79 => x"23248101",
          80 => x"23261102",
          81 => x"93040500",
          82 => x"13040000",
          83 => x"130989bb",
          84 => x"930a5001",
          85 => x"938bf5ff",
          86 => x"130bf007",
          87 => x"130a2000",
          88 => x"93092001",
          89 => x"371c0010",
          90 => x"eff01ff9",
          91 => x"1377f50f",
          92 => x"63c4ea0a",
          93 => x"6354ea04",
          94 => x"9307d7ff",
          95 => x"63e0f904",
          96 => x"93972700",
          97 => x"b307f900",
          98 => x"83a70700",
          99 => x"67800700",
         100 => x"630a0400",
         101 => x"1304f4ff",
         102 => x"1305f007",
         103 => x"ef000013",
         104 => x"e31a04fe",
         105 => x"eff05ff5",
         106 => x"1377f50f",
         107 => x"13040000",
         108 => x"e3d2eafc",
         109 => x"9307f007",
         110 => x"630ef70c",
         111 => x"63547405",
         112 => x"9377f50f",
         113 => x"938607fe",
         114 => x"93f6f60f",
         115 => x"1306e005",
         116 => x"e36cd6f8",
         117 => x"b3868400",
         118 => x"13050700",
         119 => x"2380f600",
         120 => x"ef00c00e",
         121 => x"eff05ff1",
         122 => x"1377f50f",
         123 => x"93075001",
         124 => x"13041400",
         125 => x"e3d0e7f8",
         126 => x"9307f007",
         127 => x"6302f702",
         128 => x"e34074fd",
         129 => x"13057000",
         130 => x"ef00400c",
         131 => x"eff0dfee",
         132 => x"1377f50f",
         133 => x"e3d0eaf6",
         134 => x"e31267fb",
         135 => x"630c0406",
         136 => x"1305f007",
         137 => x"ef00800a",
         138 => x"1304f4ff",
         139 => x"6ff0dff3",
         140 => x"b3848400",
         141 => x"37150010",
         142 => x"23800400",
         143 => x"130545c2",
         144 => x"ef00c00a",
         145 => x"8320c102",
         146 => x"13050400",
         147 => x"03248102",
         148 => x"83244102",
         149 => x"03290102",
         150 => x"8329c101",
         151 => x"032a8101",
         152 => x"832a4101",
         153 => x"032b0101",
         154 => x"832bc100",
         155 => x"032c8100",
         156 => x"13010103",
         157 => x"67800000",
         158 => x"1305ccf0",
         159 => x"ef000007",
         160 => x"eff09fe7",
         161 => x"1377f50f",
         162 => x"13040000",
         163 => x"e3d4eaee",
         164 => x"6ff05ff2",
         165 => x"13057000",
         166 => x"ef004003",
         167 => x"6ff09ff0",
         168 => x"f32710fc",
         169 => x"63960700",
         170 => x"b7f7fa02",
         171 => x"93870708",
         172 => x"63060500",
         173 => x"33d5a702",
         174 => x"1305f5ff",
         175 => x"b70700f0",
         176 => x"23a6a702",
         177 => x"23a0b702",
         178 => x"67800000",
         179 => x"1375f50f",
         180 => x"b70700f0",
         181 => x"370700f0",
         182 => x"23a4a702",
         183 => x"83274702",
         184 => x"93f70701",
         185 => x"e38c07fe",
         186 => x"67800000",
         187 => x"630e0502",
         188 => x"130101ff",
         189 => x"23248100",
         190 => x"23261100",
         191 => x"13040500",
         192 => x"03450500",
         193 => x"630a0500",
         194 => x"13041400",
         195 => x"eff01ffc",
         196 => x"03450400",
         197 => x"e31a05fe",
         198 => x"8320c100",
         199 => x"03248100",
         200 => x"13010101",
         201 => x"67800000",
         202 => x"67800000",
         203 => x"130101fe",
         204 => x"232e1100",
         205 => x"232c8100",
         206 => x"232a9100",
         207 => x"23282101",
         208 => x"23263101",
         209 => x"23244101",
         210 => x"6358a008",
         211 => x"b7190010",
         212 => x"13090500",
         213 => x"93040000",
         214 => x"13040000",
         215 => x"938999e0",
         216 => x"130a1000",
         217 => x"6f000001",
         218 => x"3364c400",
         219 => x"93841400",
         220 => x"63029904",
         221 => x"eff05fd8",
         222 => x"b387a900",
         223 => x"83c70700",
         224 => x"130605fd",
         225 => x"13144400",
         226 => x"13f74700",
         227 => x"93f64704",
         228 => x"e31c07fc",
         229 => x"93f73700",
         230 => x"e38a06fc",
         231 => x"63944701",
         232 => x"13050502",
         233 => x"130595fa",
         234 => x"93841400",
         235 => x"3364a400",
         236 => x"e31299fc",
         237 => x"8320c101",
         238 => x"13050400",
         239 => x"03248101",
         240 => x"83244101",
         241 => x"03290101",
         242 => x"8329c100",
         243 => x"032a8100",
         244 => x"13010102",
         245 => x"67800000",
         246 => x"13040000",
         247 => x"6ff09ffd",
         248 => x"83470500",
         249 => x"37160010",
         250 => x"130696e0",
         251 => x"3307f600",
         252 => x"03470700",
         253 => x"93060500",
         254 => x"13758700",
         255 => x"630e0500",
         256 => x"83c71600",
         257 => x"93861600",
         258 => x"3307f600",
         259 => x"03470700",
         260 => x"13758700",
         261 => x"e31605fe",
         262 => x"13754704",
         263 => x"630a0506",
         264 => x"13050000",
         265 => x"13031000",
         266 => x"6f000002",
         267 => x"83c71600",
         268 => x"33e5a800",
         269 => x"93861600",
         270 => x"3307f600",
         271 => x"03470700",
         272 => x"13784704",
         273 => x"63000804",
         274 => x"13784700",
         275 => x"938807fd",
         276 => x"13773700",
         277 => x"13154500",
         278 => x"e31a08fc",
         279 => x"63146700",
         280 => x"93870702",
         281 => x"938797fa",
         282 => x"33e5a700",
         283 => x"83c71600",
         284 => x"93861600",
         285 => x"3307f600",
         286 => x"03470700",
         287 => x"13784704",
         288 => x"e31408fc",
         289 => x"63840500",
         290 => x"23a0d500",
         291 => x"67800000",
         292 => x"13050000",
         293 => x"6ff01fff",
         294 => x"130101fe",
         295 => x"232e1100",
         296 => x"232c8100",
         297 => x"23220100",
         298 => x"23240100",
         299 => x"23260100",
         300 => x"63000506",
         301 => x"13040500",
         302 => x"63440504",
         303 => x"93074100",
         304 => x"9306a000",
         305 => x"93059000",
         306 => x"3377d402",
         307 => x"13850700",
         308 => x"9387f7ff",
         309 => x"13060400",
         310 => x"13070703",
         311 => x"a385e700",
         312 => x"3354d402",
         313 => x"e3e2c5fe",
         314 => x"3305d500",
         315 => x"eff01fe0",
         316 => x"8320c101",
         317 => x"03248101",
         318 => x"13010102",
         319 => x"67800000",
         320 => x"1305d002",
         321 => x"eff09fdc",
         322 => x"33048040",
         323 => x"6ff01ffb",
         324 => x"13050003",
         325 => x"eff09fdb",
         326 => x"8320c101",
         327 => x"03248101",
         328 => x"13010102",
         329 => x"67800000",
         330 => x"130101fe",
         331 => x"232e1100",
         332 => x"23220100",
         333 => x"23240100",
         334 => x"23060100",
         335 => x"9387f5ff",
         336 => x"13077000",
         337 => x"6376f700",
         338 => x"93077000",
         339 => x"93058000",
         340 => x"13074100",
         341 => x"b307f700",
         342 => x"b385b740",
         343 => x"13069003",
         344 => x"9376f500",
         345 => x"13870603",
         346 => x"6374e600",
         347 => x"13877605",
         348 => x"2380e700",
         349 => x"9387f7ff",
         350 => x"13554500",
         351 => x"e392f5fe",
         352 => x"13054100",
         353 => x"eff09fd6",
         354 => x"8320c101",
         355 => x"13010102",
         356 => x"67800000",
         357 => x"37c50100",
         358 => x"130101f8",
         359 => x"93050000",
         360 => x"13050520",
         361 => x"232e1106",
         362 => x"232c8106",
         363 => x"232a9106",
         364 => x"23282107",
         365 => x"23263107",
         366 => x"23244107",
         367 => x"23225107",
         368 => x"23206107",
         369 => x"232e7105",
         370 => x"232c8105",
         371 => x"232a9105",
         372 => x"2328a105",
         373 => x"2326b105",
         374 => x"eff09fcc",
         375 => x"37150010",
         376 => x"130545c0",
         377 => x"eff09fd0",
         378 => x"37150010",
         379 => x"130585c2",
         380 => x"eff0dfcf",
         381 => x"732510fc",
         382 => x"37190010",
         383 => x"eff0dfe9",
         384 => x"130549c2",
         385 => x"eff09fce",
         386 => x"b70700f0",
         387 => x"1307f03f",
         388 => x"370a1000",
         389 => x"b709a000",
         390 => x"23a2e700",
         391 => x"93041000",
         392 => x"130afaff",
         393 => x"b70a00f0",
         394 => x"93891900",
         395 => x"b3f74401",
         396 => x"639c0700",
         397 => x"1305a002",
         398 => x"eff05fc9",
         399 => x"83a74a00",
         400 => x"93d71700",
         401 => x"23a2fa00",
         402 => x"eff01faa",
         403 => x"13040500",
         404 => x"631a050c",
         405 => x"93841400",
         406 => x"e39a34fd",
         407 => x"b70700f0",
         408 => x"23a20700",
         409 => x"631a0400",
         410 => x"93050000",
         411 => x"13050000",
         412 => x"eff01fc3",
         413 => x"e7000400",
         414 => x"eff01fa8",
         415 => x"93071002",
         416 => x"93040000",
         417 => x"631cf51c",
         418 => x"37140010",
         419 => x"1305c4c3",
         420 => x"eff0dfc5",
         421 => x"b70900f0",
         422 => x"930a3005",
         423 => x"130ba004",
         424 => x"930b3002",
         425 => x"130a2000",
         426 => x"130ca000",
         427 => x"83a74900",
         428 => x"93c71700",
         429 => x"23a2f900",
         430 => x"eff01fa4",
         431 => x"1375f50f",
         432 => x"63185517",
         433 => x"eff05fa3",
         434 => x"937cf50f",
         435 => x"9387fcfc",
         436 => x"93f7f70f",
         437 => x"6360fa10",
         438 => x"93071003",
         439 => x"6398fc04",
         440 => x"13052000",
         441 => x"eff09fc4",
         442 => x"130dd5ff",
         443 => x"13054000",
         444 => x"eff0dfc3",
         445 => x"b70d01ff",
         446 => x"930c0500",
         447 => x"330dad00",
         448 => x"938dfdff",
         449 => x"639aac05",
         450 => x"930ca000",
         451 => x"eff0df9e",
         452 => x"1375f50f",
         453 => x"e31c95ff",
         454 => x"1305c4c3",
         455 => x"eff01fbd",
         456 => x"6ff0dff8",
         457 => x"13041000",
         458 => x"6ff05ff3",
         459 => x"93072003",
         460 => x"13052000",
         461 => x"639afc00",
         462 => x"eff05fbf",
         463 => x"130dc5ff",
         464 => x"13056000",
         465 => x"6ff0dffa",
         466 => x"eff05fbe",
         467 => x"130db5ff",
         468 => x"13058000",
         469 => x"6ff0dff9",
         470 => x"93f5ccff",
         471 => x"13052000",
         472 => x"2326b100",
         473 => x"eff09fbc",
         474 => x"8325c100",
         475 => x"93070500",
         476 => x"b7060001",
         477 => x"3706ffff",
         478 => x"13f53c00",
         479 => x"03a70500",
         480 => x"13083000",
         481 => x"9386f6ff",
         482 => x"93081000",
         483 => x"1306f60f",
         484 => x"63064503",
         485 => x"630a0503",
         486 => x"630c1501",
         487 => x"137707f0",
         488 => x"b3e7e700",
         489 => x"23a0f500",
         490 => x"938c1c00",
         491 => x"6ff09ff5",
         492 => x"3377c700",
         493 => x"93978700",
         494 => x"6ff09ffe",
         495 => x"3377b701",
         496 => x"93970701",
         497 => x"6ff0dffd",
         498 => x"3377d700",
         499 => x"93978701",
         500 => x"6ff01ffd",
         501 => x"93879cfc",
         502 => x"93f7f70f",
         503 => x"6362fa04",
         504 => x"13052000",
         505 => x"eff09fb4",
         506 => x"93077003",
         507 => x"13058000",
         508 => x"638afc00",
         509 => x"93078003",
         510 => x"13056000",
         511 => x"6384fc00",
         512 => x"13054000",
         513 => x"eff09fb2",
         514 => x"93040500",
         515 => x"930ca000",
         516 => x"eff09f8e",
         517 => x"1375f50f",
         518 => x"e31c95ff",
         519 => x"6ff0dfef",
         520 => x"eff09f8d",
         521 => x"1375f50f",
         522 => x"e31c85ff",
         523 => x"6ff0dfee",
         524 => x"63186509",
         525 => x"1305c4c3",
         526 => x"eff05fab",
         527 => x"93050000",
         528 => x"13050000",
         529 => x"eff0dfa5",
         530 => x"23a20900",
         531 => x"e7800400",
         532 => x"b70700f0",
         533 => x"1307a00a",
         534 => x"23a2e700",
         535 => x"130549c2",
         536 => x"b7190010",
         537 => x"eff09fa8",
         538 => x"13040000",
         539 => x"371b0010",
         540 => x"b71b0010",
         541 => x"938999e0",
         542 => x"b7170010",
         543 => x"138507c4",
         544 => x"eff0dfa6",
         545 => x"93059002",
         546 => x"13054101",
         547 => x"eff09f88",
         548 => x"13054101",
         549 => x"ef00c02c",
         550 => x"b7170010",
         551 => x"130a0500",
         552 => x"938547c4",
         553 => x"13054101",
         554 => x"eff0df81",
         555 => x"631e0500",
         556 => x"37150010",
         557 => x"130585c4",
         558 => x"eff05fa3",
         559 => x"6f004003",
         560 => x"e31c75e5",
         561 => x"6ff0dff8",
         562 => x"b7170010",
         563 => x"938547d3",
         564 => x"13054101",
         565 => x"eff00fff",
         566 => x"63100502",
         567 => x"93050000",
         568 => x"eff01f9c",
         569 => x"b70700f0",
         570 => x"23a20700",
         571 => x"e7800400",
         572 => x"e3040af8",
         573 => x"6f004018",
         574 => x"b7170010",
         575 => x"13063000",
         576 => x"938587d3",
         577 => x"13054101",
         578 => x"ef004027",
         579 => x"63100504",
         580 => x"93050000",
         581 => x"13057101",
         582 => x"eff09fac",
         583 => x"93773500",
         584 => x"13040500",
         585 => x"63940706",
         586 => x"93058000",
         587 => x"eff0dfbf",
         588 => x"37150010",
         589 => x"1305c5d3",
         590 => x"eff05f9b",
         591 => x"03250400",
         592 => x"93058000",
         593 => x"eff05fbe",
         594 => x"6ff09ffa",
         595 => x"13063000",
         596 => x"93058bd5",
         597 => x"13054101",
         598 => x"ef004022",
         599 => x"631e0502",
         600 => x"93050101",
         601 => x"13057101",
         602 => x"eff09fa7",
         603 => x"93773500",
         604 => x"13040500",
         605 => x"639c0700",
         606 => x"03250101",
         607 => x"93050000",
         608 => x"eff01fa6",
         609 => x"2320a400",
         610 => x"6ff09ff6",
         611 => x"37150010",
         612 => x"130505d4",
         613 => x"6ff05ff2",
         614 => x"13063000",
         615 => x"9385cbd5",
         616 => x"13054101",
         617 => x"ef00801d",
         618 => x"83474101",
         619 => x"1307e006",
         620 => x"630c0508",
         621 => x"639ae70a",
         622 => x"93773400",
         623 => x"e39807fc",
         624 => x"130c0404",
         625 => x"b71c0010",
         626 => x"371d0010",
         627 => x"930d80ff",
         628 => x"93058000",
         629 => x"13050400",
         630 => x"eff01fb5",
         631 => x"1385ccd3",
         632 => x"eff0df90",
         633 => x"83270400",
         634 => x"93058000",
         635 => x"130a8001",
         636 => x"13850700",
         637 => x"2326f100",
         638 => x"eff01fb3",
         639 => x"13050dd6",
         640 => x"eff0df8e",
         641 => x"b70a00ff",
         642 => x"8327c100",
         643 => x"33f55701",
         644 => x"33554501",
         645 => x"b3063501",
         646 => x"83c60600",
         647 => x"93f67609",
         648 => x"63800604",
         649 => x"130a8aff",
         650 => x"eff05f8a",
         651 => x"93da8a00",
         652 => x"e31cbafd",
         653 => x"13044400",
         654 => x"130549c2",
         655 => x"eff01f8b",
         656 => x"e31884f9",
         657 => x"6ff05fe3",
         658 => x"e388e7f6",
         659 => x"93050000",
         660 => x"13057101",
         661 => x"eff0df98",
         662 => x"13040500",
         663 => x"6ff0dff5",
         664 => x"1305e002",
         665 => x"6ff01ffc",
         666 => x"e3080ae0",
         667 => x"37150010",
         668 => x"130545d6",
         669 => x"eff09f87",
         670 => x"130549c2",
         671 => x"eff01f87",
         672 => x"6ff09fdf",
         673 => x"130101ff",
         674 => x"23248100",
         675 => x"23261100",
         676 => x"93070000",
         677 => x"13040500",
         678 => x"63880700",
         679 => x"93050000",
         680 => x"97000000",
         681 => x"e7000000",
         682 => x"b7170010",
         683 => x"03a587f1",
         684 => x"83278502",
         685 => x"63840700",
         686 => x"e7800700",
         687 => x"13050400",
         688 => x"eff04fe2",
         689 => x"130101ff",
         690 => x"23248100",
         691 => x"23229100",
         692 => x"37140010",
         693 => x"b7140010",
         694 => x"9387c4f1",
         695 => x"1304c4f1",
         696 => x"3304f440",
         697 => x"23202101",
         698 => x"23261100",
         699 => x"13542440",
         700 => x"9384c4f1",
         701 => x"13090000",
         702 => x"63108904",
         703 => x"b7140010",
         704 => x"37140010",
         705 => x"9387c4f1",
         706 => x"1304c4f1",
         707 => x"3304f440",
         708 => x"13542440",
         709 => x"9384c4f1",
         710 => x"13090000",
         711 => x"63188902",
         712 => x"8320c100",
         713 => x"03248100",
         714 => x"83244100",
         715 => x"03290100",
         716 => x"13010101",
         717 => x"67800000",
         718 => x"83a70400",
         719 => x"13091900",
         720 => x"93844400",
         721 => x"e7800700",
         722 => x"6ff01ffb",
         723 => x"83a70400",
         724 => x"13091900",
         725 => x"93844400",
         726 => x"e7800700",
         727 => x"6ff01ffc",
         728 => x"93070500",
         729 => x"03c70700",
         730 => x"93871700",
         731 => x"e31c07fe",
         732 => x"3385a740",
         733 => x"1305f5ff",
         734 => x"67800000",
         735 => x"630a0602",
         736 => x"1306f6ff",
         737 => x"13070000",
         738 => x"b307e500",
         739 => x"b386e500",
         740 => x"83c70700",
         741 => x"83c60600",
         742 => x"6398d700",
         743 => x"6306c700",
         744 => x"13071700",
         745 => x"e39207fe",
         746 => x"3385d740",
         747 => x"67800000",
         748 => x"13050000",
         749 => x"67800000",
         750 => x"78020010",
         751 => x"bc010010",
         752 => x"bc010010",
         753 => x"bc010010",
         754 => x"bc010010",
         755 => x"1c020010",
         756 => x"bc010010",
         757 => x"30020010",
         758 => x"bc010010",
         759 => x"bc010010",
         760 => x"30020010",
         761 => x"bc010010",
         762 => x"bc010010",
         763 => x"bc010010",
         764 => x"bc010010",
         765 => x"bc010010",
         766 => x"bc010010",
         767 => x"bc010010",
         768 => x"90010010",
         769 => x"0d0a5448",
         770 => x"55415320",
         771 => x"52495343",
         772 => x"2d562042",
         773 => x"6f6f746c",
         774 => x"6f616465",
         775 => x"72207630",
         776 => x"2e342e31",
         777 => x"0d0a0000",
         778 => x"436c6f63",
         779 => x"6b206672",
         780 => x"65717565",
         781 => x"6e63793a",
         782 => x"20000000",
         783 => x"3f0a0000",
         784 => x"3e200000",
         785 => x"68000000",
         786 => x"48656c70",
         787 => x"3a0d0a20",
         788 => x"68202020",
         789 => x"20202020",
         790 => x"20202020",
         791 => x"20202020",
         792 => x"202d2074",
         793 => x"68697320",
         794 => x"68656c70",
         795 => x"0d0a2072",
         796 => x"20202020",
         797 => x"20202020",
         798 => x"20202020",
         799 => x"20202020",
         800 => x"2d207275",
         801 => x"6e206170",
         802 => x"706c6963",
         803 => x"6174696f",
         804 => x"6e0d0a20",
         805 => x"7277203c",
         806 => x"61646472",
         807 => x"3e202020",
         808 => x"20202020",
         809 => x"202d2072",
         810 => x"65616420",
         811 => x"776f7264",
         812 => x"2066726f",
         813 => x"6d206164",
         814 => x"64720d0a",
         815 => x"20777720",
         816 => x"3c616464",
         817 => x"723e203c",
         818 => x"64617461",
         819 => x"3e202d20",
         820 => x"77726974",
         821 => x"6520776f",
         822 => x"72642064",
         823 => x"61746120",
         824 => x"61742061",
         825 => x"6464720d",
         826 => x"0a206477",
         827 => x"203c6164",
         828 => x"64723e20",
         829 => x"20202020",
         830 => x"2020202d",
         831 => x"2064756d",
         832 => x"70203136",
         833 => x"20776f72",
         834 => x"64730d0a",
         835 => x"206e2020",
         836 => x"20202020",
         837 => x"20202020",
         838 => x"20202020",
         839 => x"20202d20",
         840 => x"64756d70",
         841 => x"206e6578",
         842 => x"74203136",
         843 => x"20776f72",
         844 => x"64730000",
         845 => x"72000000",
         846 => x"72772000",
         847 => x"3a200000",
         848 => x"4e6f7420",
         849 => x"6f6e2034",
         850 => x"2d627974",
         851 => x"6520626f",
         852 => x"756e6461",
         853 => x"72792100",
         854 => x"77772000",
         855 => x"64772000",
         856 => x"20200000",
         857 => x"3f3f0000",
         858 => x"626f6f74",
         859 => x"6c6f6164",
         860 => x"65720000",
         861 => x"54485541",
         862 => x"53205249",
         863 => x"53432d56",
         864 => x"20525633",
         865 => x"32494d20",
         866 => x"62617265",
         867 => x"206d6574",
         868 => x"616c2070",
         869 => x"726f6365",
         870 => x"73736f72",
         871 => x"00000000",
         872 => x"54686520",
         873 => x"48616775",
         874 => x"6520556e",
         875 => x"69766572",
         876 => x"73697479",
         877 => x"206f6620",
         878 => x"4170706c",
         879 => x"69656420",
         880 => x"53636965",
         881 => x"6e636573",
         882 => x"00000000",
         883 => x"44657061",
         884 => x"72746d65",
         885 => x"6e74206f",
         886 => x"6620456c",
         887 => x"65637472",
         888 => x"6963616c",
         889 => x"20456e67",
         890 => x"696e6565",
         891 => x"72696e67",
         892 => x"00000000",
         893 => x"4a2e452e",
         894 => x"4a2e206f",
         895 => x"70206465",
         896 => x"6e204272",
         897 => x"6f757700",
         898 => x"00202020",
         899 => x"20202020",
         900 => x"20202828",
         901 => x"28282820",
         902 => x"20202020",
         903 => x"20202020",
         904 => x"20202020",
         905 => x"20202020",
         906 => x"20881010",
         907 => x"10101010",
         908 => x"10101010",
         909 => x"10101010",
         910 => x"10040404",
         911 => x"04040404",
         912 => x"04040410",
         913 => x"10101010",
         914 => x"10104141",
         915 => x"41414141",
         916 => x"01010101",
         917 => x"01010101",
         918 => x"01010101",
         919 => x"01010101",
         920 => x"01010101",
         921 => x"10101010",
         922 => x"10104242",
         923 => x"42424242",
         924 => x"02020202",
         925 => x"02020202",
         926 => x"02020202",
         927 => x"02020202",
         928 => x"02020202",
         929 => x"10101010",
         930 => x"20000000",
         931 => x"00000000",
         932 => x"00000000",
         933 => x"00000000",
         934 => x"00000000",
         935 => x"00000000",
         936 => x"00000000",
         937 => x"00000000",
         938 => x"00000000",
         939 => x"00000000",
         940 => x"00000000",
         941 => x"00000000",
         942 => x"00000000",
         943 => x"00000000",
         944 => x"00000000",
         945 => x"00000000",
         946 => x"00000000",
         947 => x"00000000",
         948 => x"00000000",
         949 => x"00000000",
         950 => x"00000000",
         951 => x"00000000",
         952 => x"00000000",
         953 => x"00000000",
         954 => x"00000000",
         955 => x"00000000",
         956 => x"00000000",
         957 => x"00000000",
         958 => x"00000000",
         959 => x"00000000",
         960 => x"00000000",
         961 => x"00000000",
         962 => x"00000000",
         963 => x"3c627265",
         964 => x"616b3e0d",
         965 => x"0a000000",
         966 => x"18000020",
         967 => x"680d0010",
         968 => x"740d0010",
         969 => x"a00d0010",
         970 => x"cc0d0010",
         971 => x"f40d0010",
         972 => x"00000000",
         973 => x"00000000",
         974 => x"00000000",
         975 => x"00000000",
         976 => x"00000000",
         977 => x"00000000",
         978 => x"00000000",
         979 => x"00000000",
         980 => x"00000000",
         981 => x"00000000",
         982 => x"00000000",
         983 => x"00000000",
         984 => x"00000000",
         985 => x"00000000",
         986 => x"00000000",
         987 => x"00000000",
         988 => x"00000000",
         989 => x"00000000",
         990 => x"00000000",
         991 => x"00000000",
         992 => x"00000000",
         993 => x"00000000",
         994 => x"00000000",
         995 => x"00000000",
         996 => x"00000000",
         997 => x"18000020",
         others => (others => '0')
        );

begin

    gen_bootrom: if HAVE_BOOTLOADER_ROM generate

        -- ROM, for both instructions and read-only data
        process (I_clk, I_areset, I_pc, I_memaddress, I_csboot, I_memsize, I_stall) is
        variable address_instr : integer range 0 to bootloader_size-1;
        variable address_data : integer range 0 to bootloader_size-1;
        variable instr_var : data_type;
        variable instr_recode : data_type;
        variable romdata_var : data_type;
        constant x : data_type := (others => 'X');
        begin
            -- Calculate addresses
            address_instr := to_integer(unsigned(I_pc(bootloader_size_bits-1 downto 2)));
            address_data := to_integer(unsigned(I_memaddress(bootloader_size_bits-1 downto 2)));

            -- Quartus will detect ROM table and uses onboard RAM
            -- Do not use reset, otherwise ROM will be created with ALMs
            if rising_edge(I_clk) then
                if I_stall = '0' then
                    instr_var := bootrom(address_instr);
                end if;
                romdata_var := bootrom(address_data);
            end if;
            
            -- Recode instruction
            O_instr <= instr_var(7 downto 0) & instr_var(15 downto 8) & instr_var(23 downto 16) & instr_var(31 downto 24);
            
            O_load_misaligned_error <= '0';
            
            -- By natural size, for data
            if I_csboot = '1' then
                if I_memsize = memsize_word and I_memaddress(1 downto 0) = "00" then
                    O_dataout <= romdata_var(7 downto 0) & romdata_var(15 downto 8) & romdata_var(23 downto 16) & romdata_var(31 downto 24);
                elsif I_memsize = memsize_halfword and I_memaddress(1 downto 0) = "00" then
                    O_dataout <= x(31 downto 16) & romdata_var(23 downto 16) & romdata_var(31 downto 24);
                elsif I_memsize = memsize_halfword and I_memaddress(1 downto 0) = "10" then
                    O_dataout <= x(31 downto 16) & romdata_var(7 downto 0) & romdata_var(15 downto 8);
                elsif I_memsize = memsize_byte then
                    case I_memaddress(1 downto 0) is
                        when "00" => O_dataout <= x(31 downto 8) & romdata_var(31 downto 24);
                        when "01" => O_dataout <= x(31 downto 8) & romdata_var(23 downto 16);
                        when "10" => O_dataout <= x(31 downto 8) & romdata_var(15 downto 8);
                        when "11" => O_dataout <= x(31 downto 8) & romdata_var(7 downto 0);
                        when others => O_dataout <= x; O_load_misaligned_error <= '1';
                    end case;
                else
                    -- Chip select, but not aligned
                    O_dataout <= x;
                    O_load_misaligned_error <= '1';
                end if;
            else
                -- No chip select, so no data
                O_dataout <= x;
            end if;
        end process;
    end generate;

    gen_bootrom_not: if not HAVE_BOOTLOADER_ROM generate
        O_load_misaligned_error <= '0';
        O_dataout <= (others => 'X');
        O_instr  <= (others => 'X');
    end generate;
end architecture rtl;
