-- srec2vhdl table generator
-- for input file interrupt_direct.srec

library ieee;
use ieee.std_logic_1164.all;

library work;
use work.processor_common.all;

package processor_common_rom is
    constant rom_contents : rom_type := (
           0 => x"97020000",
           1 => x"93828226",
           2 => x"73905230",
           3 => x"97010020",
           4 => x"9381417f",
           5 => x"17810020",
           6 => x"1301c1fe",
           7 => x"13860188",
           8 => x"93874189",
           9 => x"637af600",
          10 => x"3386c740",
          11 => x"93050000",
          12 => x"13850188",
          13 => x"ef10002f",
          14 => x"37050020",
          15 => x"13060500",
          16 => x"93870188",
          17 => x"637cf600",
          18 => x"b7350000",
          19 => x"3386c740",
          20 => x"9385c5fe",
          21 => x"13050500",
          22 => x"ef10802a",
          23 => x"ef10c07e",
          24 => x"b7050020",
          25 => x"13060000",
          26 => x"93850500",
          27 => x"13055000",
          28 => x"ef100049",
          29 => x"ef104079",
          30 => x"6f10c03f",
          31 => x"130101ff",
          32 => x"23261100",
          33 => x"ef10c041",
          34 => x"8320c100",
          35 => x"13051000",
          36 => x"13010101",
          37 => x"67800000",
          38 => x"130101fd",
          39 => x"232c4101",
          40 => x"130a0500",
          41 => x"37350000",
          42 => x"130585e3",
          43 => x"23248102",
          44 => x"23229102",
          45 => x"23202103",
          46 => x"232e3101",
          47 => x"83244a08",
          48 => x"23261102",
          49 => x"13044100",
          50 => x"ef10803f",
          51 => x"37390000",
          52 => x"9309c1ff",
          53 => x"93070400",
          54 => x"1309c9c0",
          55 => x"13f7f400",
          56 => x"3307e900",
          57 => x"03470700",
          58 => x"9387f7ff",
          59 => x"93d44400",
          60 => x"2384e700",
          61 => x"e39437ff",
          62 => x"13054100",
          63 => x"23060100",
          64 => x"ef10003c",
          65 => x"37350000",
          66 => x"1305c5e4",
          67 => x"ef10403b",
          68 => x"03278a08",
          69 => x"9377f700",
          70 => x"b307f900",
          71 => x"83c70700",
          72 => x"1304f4ff",
          73 => x"13574700",
          74 => x"2304f400",
          75 => x"e31434ff",
          76 => x"13054100",
          77 => x"ef10c038",
          78 => x"37350000",
          79 => x"130545e8",
          80 => x"ef100038",
          81 => x"8320c102",
          82 => x"03248102",
          83 => x"83244102",
          84 => x"03290102",
          85 => x"8329c101",
          86 => x"032a8101",
          87 => x"13010103",
          88 => x"67800000",
          89 => x"b70700f0",
          90 => x"03a74708",
          91 => x"1377f7fe",
          92 => x"23a2e708",
          93 => x"03a74700",
          94 => x"13471700",
          95 => x"23a2e700",
          96 => x"67800000",
          97 => x"370700f0",
          98 => x"83274700",
          99 => x"93e70720",
         100 => x"2322f700",
         101 => x"6f000000",
         102 => x"b70700f0",
         103 => x"83a6470f",
         104 => x"03a6070f",
         105 => x"03a7470f",
         106 => x"e31ad7fe",
         107 => x"b7860100",
         108 => x"9305f0ff",
         109 => x"9386066a",
         110 => x"23aeb70e",
         111 => x"b306d600",
         112 => x"23acb70e",
         113 => x"33b6c600",
         114 => x"23acd70e",
         115 => x"3306e600",
         116 => x"23aec70e",
         117 => x"03a74700",
         118 => x"13472700",
         119 => x"23a2e700",
         120 => x"67800000",
         121 => x"b70700f0",
         122 => x"03a74702",
         123 => x"13774700",
         124 => x"630a0700",
         125 => x"03a74700",
         126 => x"13478700",
         127 => x"23a2e700",
         128 => x"83a78702",
         129 => x"67800000",
         130 => x"b70700f0",
         131 => x"03a7470a",
         132 => x"1377f7f0",
         133 => x"23a2e70a",
         134 => x"03a74700",
         135 => x"13474700",
         136 => x"23a2e700",
         137 => x"67800000",
         138 => x"b70700f0",
         139 => x"03a74706",
         140 => x"137777ff",
         141 => x"23a2e706",
         142 => x"03a74700",
         143 => x"13470701",
         144 => x"23a2e700",
         145 => x"67800000",
         146 => x"b70700f0",
         147 => x"03a74704",
         148 => x"137777fe",
         149 => x"23a2e704",
         150 => x"03a74700",
         151 => x"13470702",
         152 => x"23a2e700",
         153 => x"67800000",
         154 => x"6f000000",
         155 => x"13050000",
         156 => x"67800000",
         157 => x"13050000",
         158 => x"67800000",
         159 => x"130101f7",
         160 => x"23221100",
         161 => x"23242100",
         162 => x"23263100",
         163 => x"23284100",
         164 => x"232a5100",
         165 => x"232c6100",
         166 => x"232e7100",
         167 => x"23208102",
         168 => x"23229102",
         169 => x"2324a102",
         170 => x"2326b102",
         171 => x"2328c102",
         172 => x"232ad102",
         173 => x"232ce102",
         174 => x"232ef102",
         175 => x"23200105",
         176 => x"23221105",
         177 => x"23242105",
         178 => x"23263105",
         179 => x"23284105",
         180 => x"232a5105",
         181 => x"232c6105",
         182 => x"232e7105",
         183 => x"23208107",
         184 => x"23229107",
         185 => x"2324a107",
         186 => x"2326b107",
         187 => x"2328c107",
         188 => x"232ad107",
         189 => x"232ce107",
         190 => x"232ef107",
         191 => x"f3222034",
         192 => x"23205108",
         193 => x"f3221034",
         194 => x"23225108",
         195 => x"83a20200",
         196 => x"23245108",
         197 => x"f3223034",
         198 => x"23265108",
         199 => x"f3272034",
         200 => x"37070080",
         201 => x"93067700",
         202 => x"6380d710",
         203 => x"9306b000",
         204 => x"63fef602",
         205 => x"934607ff",
         206 => x"b386d700",
         207 => x"13065000",
         208 => x"636ad602",
         209 => x"1347f7fe",
         210 => x"b387e700",
         211 => x"13074000",
         212 => x"6364f716",
         213 => x"37370000",
         214 => x"93972700",
         215 => x"130707c2",
         216 => x"b387e700",
         217 => x"83a70700",
         218 => x"67800700",
         219 => x"13071000",
         220 => x"636ef708",
         221 => x"03258102",
         222 => x"83220108",
         223 => x"63c80200",
         224 => x"f3221034",
         225 => x"93824200",
         226 => x"73901234",
         227 => x"832fc107",
         228 => x"032f8107",
         229 => x"832e4107",
         230 => x"032e0107",
         231 => x"832dc106",
         232 => x"032d8106",
         233 => x"832c4106",
         234 => x"032c0106",
         235 => x"832bc105",
         236 => x"032b8105",
         237 => x"832a4105",
         238 => x"032a0105",
         239 => x"8329c104",
         240 => x"03298104",
         241 => x"83284104",
         242 => x"03280104",
         243 => x"8327c103",
         244 => x"03278103",
         245 => x"83264103",
         246 => x"03260103",
         247 => x"8325c102",
         248 => x"83244102",
         249 => x"03240102",
         250 => x"8323c101",
         251 => x"03238101",
         252 => x"83224101",
         253 => x"03220101",
         254 => x"8321c100",
         255 => x"03218100",
         256 => x"83204100",
         257 => x"13010109",
         258 => x"73002030",
         259 => x"e3e4f6f6",
         260 => x"37370000",
         261 => x"93972700",
         262 => x"130747c3",
         263 => x"b387e700",
         264 => x"83a70700",
         265 => x"67800700",
         266 => x"eff01fd7",
         267 => x"03258102",
         268 => x"6ff09ff4",
         269 => x"eff05fdd",
         270 => x"03258102",
         271 => x"6ff0dff3",
         272 => x"eff09fde",
         273 => x"03258102",
         274 => x"6ff01ff3",
         275 => x"eff0dfdf",
         276 => x"03258102",
         277 => x"6ff05ff2",
         278 => x"eff0dfd0",
         279 => x"03258102",
         280 => x"6ff09ff1",
         281 => x"eff01fd8",
         282 => x"03258102",
         283 => x"6ff0dff0",
         284 => x"9307600d",
         285 => x"6384f806",
         286 => x"9307900a",
         287 => x"6388f818",
         288 => x"63ca170f",
         289 => x"938878fc",
         290 => x"93074002",
         291 => x"63ec1703",
         292 => x"b7370000",
         293 => x"938747c6",
         294 => x"93982800",
         295 => x"b388f800",
         296 => x"83a70800",
         297 => x"67800700",
         298 => x"13050100",
         299 => x"eff0dfbe",
         300 => x"03258102",
         301 => x"6ff05fec",
         302 => x"eff0dfcc",
         303 => x"03258102",
         304 => x"6ff09feb",
         305 => x"ef10c033",
         306 => x"93078005",
         307 => x"2320f500",
         308 => x"9307f0ff",
         309 => x"13850700",
         310 => x"6ff01fea",
         311 => x"63120510",
         312 => x"13858189",
         313 => x"13050500",
         314 => x"6ff01fe9",
         315 => x"b7270000",
         316 => x"23a2f500",
         317 => x"93070000",
         318 => x"13850700",
         319 => x"6ff0dfe7",
         320 => x"93070000",
         321 => x"13850700",
         322 => x"6ff01fe7",
         323 => x"ef10402f",
         324 => x"93079000",
         325 => x"2320f500",
         326 => x"9307f0ff",
         327 => x"13850700",
         328 => x"6ff09fe5",
         329 => x"13090600",
         330 => x"13840500",
         331 => x"635cc000",
         332 => x"b384c500",
         333 => x"03450400",
         334 => x"13041400",
         335 => x"eff01fb4",
         336 => x"e39a84fe",
         337 => x"13050900",
         338 => x"6ff01fe3",
         339 => x"13090600",
         340 => x"13840500",
         341 => x"e358c0fe",
         342 => x"b384c500",
         343 => x"eff0dfb1",
         344 => x"2300a400",
         345 => x"13041400",
         346 => x"e31a94fe",
         347 => x"13050900",
         348 => x"6ff09fe0",
         349 => x"938808c0",
         350 => x"9307f000",
         351 => x"e3e417f5",
         352 => x"b7370000",
         353 => x"938787cf",
         354 => x"93982800",
         355 => x"b388f800",
         356 => x"83a70800",
         357 => x"67800700",
         358 => x"ef108026",
         359 => x"9307d000",
         360 => x"2320f500",
         361 => x"9307f0ff",
         362 => x"13850700",
         363 => x"6ff0dfdc",
         364 => x"ef100025",
         365 => x"93072000",
         366 => x"2320f500",
         367 => x"9307f0ff",
         368 => x"13850700",
         369 => x"6ff05fdb",
         370 => x"ef108023",
         371 => x"9307f001",
         372 => x"2320f500",
         373 => x"9307f0ff",
         374 => x"13850700",
         375 => x"6ff0dfd9",
         376 => x"b7870020",
         377 => x"93870700",
         378 => x"13070040",
         379 => x"b387e740",
         380 => x"e36af5ee",
         381 => x"ef10c020",
         382 => x"9307c000",
         383 => x"2320f500",
         384 => x"1305f0ff",
         385 => x"13050500",
         386 => x"6ff01fd7",
         387 => x"13090000",
         388 => x"93040500",
         389 => x"13040900",
         390 => x"93090900",
         391 => x"93070900",
         392 => x"732410c8",
         393 => x"f32910c0",
         394 => x"f32710c8",
         395 => x"e31af4fe",
         396 => x"37460f00",
         397 => x"13060624",
         398 => x"93060000",
         399 => x"13850900",
         400 => x"93050400",
         401 => x"ef00900d",
         402 => x"37460f00",
         403 => x"23a4a400",
         404 => x"13060624",
         405 => x"93060000",
         406 => x"13850900",
         407 => x"93050400",
         408 => x"ef00c048",
         409 => x"23a0a400",
         410 => x"23a2b400",
         411 => x"13050900",
         412 => x"6ff09fd0",
         413 => x"13030500",
         414 => x"138e0500",
         415 => x"93080000",
         416 => x"63dc0500",
         417 => x"b337a000",
         418 => x"330eb040",
         419 => x"330efe40",
         420 => x"3303a040",
         421 => x"9308f0ff",
         422 => x"63dc0600",
         423 => x"b337c000",
         424 => x"b306d040",
         425 => x"93c8f8ff",
         426 => x"b386f640",
         427 => x"3306c040",
         428 => x"13070600",
         429 => x"13080300",
         430 => x"93070e00",
         431 => x"639c0628",
         432 => x"b7350000",
         433 => x"938585d3",
         434 => x"6376ce0e",
         435 => x"b7060100",
         436 => x"6378d60c",
         437 => x"93360610",
         438 => x"93c61600",
         439 => x"93963600",
         440 => x"3355d600",
         441 => x"b385a500",
         442 => x"83c50500",
         443 => x"13050002",
         444 => x"b386d500",
         445 => x"b305d540",
         446 => x"630cd500",
         447 => x"b317be00",
         448 => x"b356d300",
         449 => x"3317b600",
         450 => x"b3e7f600",
         451 => x"3318b300",
         452 => x"93550701",
         453 => x"33deb702",
         454 => x"13160701",
         455 => x"13560601",
         456 => x"b3f7b702",
         457 => x"13050e00",
         458 => x"3303c603",
         459 => x"93960701",
         460 => x"93570801",
         461 => x"b3e7d700",
         462 => x"63fe6700",
         463 => x"b307f700",
         464 => x"1305feff",
         465 => x"63e8e700",
         466 => x"63f66700",
         467 => x"1305eeff",
         468 => x"b387e700",
         469 => x"b3876740",
         470 => x"33d3b702",
         471 => x"13180801",
         472 => x"13580801",
         473 => x"b3f7b702",
         474 => x"b3066602",
         475 => x"93970701",
         476 => x"3368f800",
         477 => x"93070300",
         478 => x"637cd800",
         479 => x"33080701",
         480 => x"9307f3ff",
         481 => x"6366e800",
         482 => x"6374d800",
         483 => x"9307e3ff",
         484 => x"13150501",
         485 => x"3365f500",
         486 => x"93050000",
         487 => x"6f00000e",
         488 => x"37050001",
         489 => x"93060001",
         490 => x"e36ca6f2",
         491 => x"93068001",
         492 => x"6ff01ff3",
         493 => x"93060000",
         494 => x"630c0600",
         495 => x"b7070100",
         496 => x"637af60c",
         497 => x"93360610",
         498 => x"93c61600",
         499 => x"93963600",
         500 => x"b357d600",
         501 => x"b385f500",
         502 => x"83c70500",
         503 => x"b387d700",
         504 => x"93060002",
         505 => x"b385f640",
         506 => x"6390f60c",
         507 => x"b307ce40",
         508 => x"93051000",
         509 => x"13530701",
         510 => x"b3de6702",
         511 => x"13160701",
         512 => x"13560601",
         513 => x"93560801",
         514 => x"b3f76702",
         515 => x"13850e00",
         516 => x"330ed603",
         517 => x"93970701",
         518 => x"b3e7f600",
         519 => x"63fec701",
         520 => x"b307f700",
         521 => x"1385feff",
         522 => x"63e8e700",
         523 => x"63f6c701",
         524 => x"1385eeff",
         525 => x"b387e700",
         526 => x"b387c741",
         527 => x"33de6702",
         528 => x"13180801",
         529 => x"13580801",
         530 => x"b3f76702",
         531 => x"b306c603",
         532 => x"93970701",
         533 => x"3368f800",
         534 => x"93070e00",
         535 => x"637cd800",
         536 => x"33080701",
         537 => x"9307feff",
         538 => x"6366e800",
         539 => x"6374d800",
         540 => x"9307eeff",
         541 => x"13150501",
         542 => x"3365f500",
         543 => x"638a0800",
         544 => x"b337a000",
         545 => x"b305b040",
         546 => x"b385f540",
         547 => x"3305a040",
         548 => x"67800000",
         549 => x"b7070001",
         550 => x"93060001",
         551 => x"e36af6f2",
         552 => x"93068001",
         553 => x"6ff0dff2",
         554 => x"3317b600",
         555 => x"b356fe00",
         556 => x"13550701",
         557 => x"331ebe00",
         558 => x"b357f300",
         559 => x"b3e7c701",
         560 => x"33dea602",
         561 => x"13160701",
         562 => x"13560601",
         563 => x"3318b300",
         564 => x"b3f6a602",
         565 => x"3303c603",
         566 => x"93950601",
         567 => x"93d60701",
         568 => x"b3e6b600",
         569 => x"93050e00",
         570 => x"63fe6600",
         571 => x"b306d700",
         572 => x"9305feff",
         573 => x"63e8e600",
         574 => x"63f66600",
         575 => x"9305eeff",
         576 => x"b386e600",
         577 => x"b3866640",
         578 => x"33d3a602",
         579 => x"93970701",
         580 => x"93d70701",
         581 => x"b3f6a602",
         582 => x"33066602",
         583 => x"93960601",
         584 => x"b3e7d700",
         585 => x"93060300",
         586 => x"63fec700",
         587 => x"b307f700",
         588 => x"9306f3ff",
         589 => x"63e8e700",
         590 => x"63f6c700",
         591 => x"9306e3ff",
         592 => x"b387e700",
         593 => x"93950501",
         594 => x"b387c740",
         595 => x"b3e5d500",
         596 => x"6ff05fea",
         597 => x"6366de18",
         598 => x"b7070100",
         599 => x"63f4f604",
         600 => x"13b70610",
         601 => x"13471700",
         602 => x"13173700",
         603 => x"b7370000",
         604 => x"b3d5e600",
         605 => x"938787d3",
         606 => x"b387b700",
         607 => x"83c70700",
         608 => x"b387e700",
         609 => x"13070002",
         610 => x"b305f740",
         611 => x"6316f702",
         612 => x"13051000",
         613 => x"e3e4c6ef",
         614 => x"3335c300",
         615 => x"13451500",
         616 => x"6ff0dfed",
         617 => x"b7070001",
         618 => x"13070001",
         619 => x"e3e0f6fc",
         620 => x"13078001",
         621 => x"6ff09ffb",
         622 => x"3357f600",
         623 => x"b396b600",
         624 => x"b366d700",
         625 => x"3357fe00",
         626 => x"331ebe00",
         627 => x"b357f300",
         628 => x"b3e7c701",
         629 => x"13de0601",
         630 => x"335fc703",
         631 => x"13980601",
         632 => x"13580801",
         633 => x"3316b600",
         634 => x"3377c703",
         635 => x"b30ee803",
         636 => x"13150701",
         637 => x"13d70701",
         638 => x"3367a700",
         639 => x"13050f00",
         640 => x"637ed701",
         641 => x"3387e600",
         642 => x"1305ffff",
         643 => x"6368d700",
         644 => x"6376d701",
         645 => x"1305efff",
         646 => x"3307d700",
         647 => x"3307d741",
         648 => x"b35ec703",
         649 => x"93970701",
         650 => x"93d70701",
         651 => x"3377c703",
         652 => x"3308d803",
         653 => x"13170701",
         654 => x"b3e7e700",
         655 => x"13870e00",
         656 => x"63fe0701",
         657 => x"b387f600",
         658 => x"1387feff",
         659 => x"63e8d700",
         660 => x"63f60701",
         661 => x"1387eeff",
         662 => x"b387d700",
         663 => x"13150501",
         664 => x"b70e0100",
         665 => x"3365e500",
         666 => x"9386feff",
         667 => x"3377d500",
         668 => x"b3870741",
         669 => x"b376d600",
         670 => x"13580501",
         671 => x"13560601",
         672 => x"330ed702",
         673 => x"b306d802",
         674 => x"3307c702",
         675 => x"3308c802",
         676 => x"3306d700",
         677 => x"13570e01",
         678 => x"3307c700",
         679 => x"6374d700",
         680 => x"3308d801",
         681 => x"93560701",
         682 => x"b3860601",
         683 => x"63e6d702",
         684 => x"e394d7ce",
         685 => x"b7070100",
         686 => x"9387f7ff",
         687 => x"3377f700",
         688 => x"13170701",
         689 => x"337efe00",
         690 => x"3313b300",
         691 => x"3307c701",
         692 => x"93050000",
         693 => x"e374e3da",
         694 => x"1305f5ff",
         695 => x"6ff0dfcb",
         696 => x"93050000",
         697 => x"13050000",
         698 => x"6ff05fd9",
         699 => x"93080500",
         700 => x"13830500",
         701 => x"13070600",
         702 => x"13080500",
         703 => x"93870500",
         704 => x"63920628",
         705 => x"b7350000",
         706 => x"938585d3",
         707 => x"6376c30e",
         708 => x"b7060100",
         709 => x"6378d60c",
         710 => x"93360610",
         711 => x"93c61600",
         712 => x"93963600",
         713 => x"3355d600",
         714 => x"b385a500",
         715 => x"83c50500",
         716 => x"13050002",
         717 => x"b386d500",
         718 => x"b305d540",
         719 => x"630cd500",
         720 => x"b317b300",
         721 => x"b3d6d800",
         722 => x"3317b600",
         723 => x"b3e7f600",
         724 => x"3398b800",
         725 => x"93550701",
         726 => x"33d3b702",
         727 => x"13160701",
         728 => x"13560601",
         729 => x"b3f7b702",
         730 => x"13050300",
         731 => x"b3086602",
         732 => x"93960701",
         733 => x"93570801",
         734 => x"b3e7d700",
         735 => x"63fe1701",
         736 => x"b307f700",
         737 => x"1305f3ff",
         738 => x"63e8e700",
         739 => x"63f61701",
         740 => x"1305e3ff",
         741 => x"b387e700",
         742 => x"b3871741",
         743 => x"b3d8b702",
         744 => x"13180801",
         745 => x"13580801",
         746 => x"b3f7b702",
         747 => x"b3061603",
         748 => x"93970701",
         749 => x"3368f800",
         750 => x"93870800",
         751 => x"637cd800",
         752 => x"33080701",
         753 => x"9387f8ff",
         754 => x"6366e800",
         755 => x"6374d800",
         756 => x"9387e8ff",
         757 => x"13150501",
         758 => x"3365f500",
         759 => x"93050000",
         760 => x"67800000",
         761 => x"37050001",
         762 => x"93060001",
         763 => x"e36ca6f2",
         764 => x"93068001",
         765 => x"6ff01ff3",
         766 => x"93060000",
         767 => x"630c0600",
         768 => x"b7070100",
         769 => x"6370f60c",
         770 => x"93360610",
         771 => x"93c61600",
         772 => x"93963600",
         773 => x"b357d600",
         774 => x"b385f500",
         775 => x"83c70500",
         776 => x"b387d700",
         777 => x"93060002",
         778 => x"b385f640",
         779 => x"6396f60a",
         780 => x"b307c340",
         781 => x"93051000",
         782 => x"93580701",
         783 => x"33de1703",
         784 => x"13160701",
         785 => x"13560601",
         786 => x"93560801",
         787 => x"b3f71703",
         788 => x"13050e00",
         789 => x"3303c603",
         790 => x"93970701",
         791 => x"b3e7f600",
         792 => x"63fe6700",
         793 => x"b307f700",
         794 => x"1305feff",
         795 => x"63e8e700",
         796 => x"63f66700",
         797 => x"1305eeff",
         798 => x"b387e700",
         799 => x"b3876740",
         800 => x"33d31703",
         801 => x"13180801",
         802 => x"13580801",
         803 => x"b3f71703",
         804 => x"b3066602",
         805 => x"93970701",
         806 => x"3368f800",
         807 => x"93070300",
         808 => x"637cd800",
         809 => x"33080701",
         810 => x"9307f3ff",
         811 => x"6366e800",
         812 => x"6374d800",
         813 => x"9307e3ff",
         814 => x"13150501",
         815 => x"3365f500",
         816 => x"67800000",
         817 => x"b7070001",
         818 => x"93060001",
         819 => x"e364f6f4",
         820 => x"93068001",
         821 => x"6ff01ff4",
         822 => x"3317b600",
         823 => x"b356f300",
         824 => x"13550701",
         825 => x"3313b300",
         826 => x"b3d7f800",
         827 => x"b3e76700",
         828 => x"33d3a602",
         829 => x"13160701",
         830 => x"13560601",
         831 => x"3398b800",
         832 => x"b3f6a602",
         833 => x"b3086602",
         834 => x"93950601",
         835 => x"93d60701",
         836 => x"b3e6b600",
         837 => x"93050300",
         838 => x"63fe1601",
         839 => x"b306d700",
         840 => x"9305f3ff",
         841 => x"63e8e600",
         842 => x"63f61601",
         843 => x"9305e3ff",
         844 => x"b386e600",
         845 => x"b3861641",
         846 => x"b3d8a602",
         847 => x"93970701",
         848 => x"93d70701",
         849 => x"b3f6a602",
         850 => x"33061603",
         851 => x"93960601",
         852 => x"b3e7d700",
         853 => x"93860800",
         854 => x"63fec700",
         855 => x"b307f700",
         856 => x"9386f8ff",
         857 => x"63e8e700",
         858 => x"63f6c700",
         859 => x"9386e8ff",
         860 => x"b387e700",
         861 => x"93950501",
         862 => x"b387c740",
         863 => x"b3e5d500",
         864 => x"6ff09feb",
         865 => x"63e6d518",
         866 => x"b7070100",
         867 => x"63f4f604",
         868 => x"13b70610",
         869 => x"13471700",
         870 => x"13173700",
         871 => x"b7370000",
         872 => x"b3d5e600",
         873 => x"938787d3",
         874 => x"b387b700",
         875 => x"83c70700",
         876 => x"b387e700",
         877 => x"13070002",
         878 => x"b305f740",
         879 => x"6316f702",
         880 => x"13051000",
         881 => x"e3ee66e0",
         882 => x"33b5c800",
         883 => x"13451500",
         884 => x"67800000",
         885 => x"b7070001",
         886 => x"13070001",
         887 => x"e3e0f6fc",
         888 => x"13078001",
         889 => x"6ff09ffb",
         890 => x"3357f600",
         891 => x"b396b600",
         892 => x"b366d700",
         893 => x"3357f300",
         894 => x"3313b300",
         895 => x"b3d7f800",
         896 => x"b3e76700",
         897 => x"13d30601",
         898 => x"b35e6702",
         899 => x"13980601",
         900 => x"13580801",
         901 => x"3316b600",
         902 => x"33776702",
         903 => x"330ed803",
         904 => x"13150701",
         905 => x"13d70701",
         906 => x"3367a700",
         907 => x"13850e00",
         908 => x"637ec701",
         909 => x"3387e600",
         910 => x"1385feff",
         911 => x"6368d700",
         912 => x"6376c701",
         913 => x"1385eeff",
         914 => x"3307d700",
         915 => x"3307c741",
         916 => x"335e6702",
         917 => x"93970701",
         918 => x"93d70701",
         919 => x"33776702",
         920 => x"3308c803",
         921 => x"13170701",
         922 => x"b3e7e700",
         923 => x"13070e00",
         924 => x"63fe0701",
         925 => x"b387f600",
         926 => x"1307feff",
         927 => x"63e8d700",
         928 => x"63f60701",
         929 => x"1307eeff",
         930 => x"b387d700",
         931 => x"13150501",
         932 => x"370e0100",
         933 => x"3365e500",
         934 => x"9306feff",
         935 => x"3377d500",
         936 => x"b3870741",
         937 => x"b376d600",
         938 => x"13580501",
         939 => x"13560601",
         940 => x"3303d702",
         941 => x"b306d802",
         942 => x"3307c702",
         943 => x"3308c802",
         944 => x"3306d700",
         945 => x"13570301",
         946 => x"3307c700",
         947 => x"6374d700",
         948 => x"3308c801",
         949 => x"93560701",
         950 => x"b3860601",
         951 => x"63e6d702",
         952 => x"e39ed7ce",
         953 => x"b7070100",
         954 => x"9387f7ff",
         955 => x"3377f700",
         956 => x"13170701",
         957 => x"3373f300",
         958 => x"b398b800",
         959 => x"33076700",
         960 => x"93050000",
         961 => x"e3fee8cc",
         962 => x"1305f5ff",
         963 => x"6ff01fcd",
         964 => x"93050000",
         965 => x"13050000",
         966 => x"67800000",
         967 => x"13080600",
         968 => x"93070500",
         969 => x"13870500",
         970 => x"63960620",
         971 => x"b7380000",
         972 => x"938888d3",
         973 => x"63fcc50c",
         974 => x"b7060100",
         975 => x"637ed60a",
         976 => x"93360610",
         977 => x"93c61600",
         978 => x"93963600",
         979 => x"3353d600",
         980 => x"b3886800",
         981 => x"83c80800",
         982 => x"13030002",
         983 => x"b386d800",
         984 => x"b308d340",
         985 => x"630cd300",
         986 => x"33971501",
         987 => x"b356d500",
         988 => x"33181601",
         989 => x"33e7e600",
         990 => x"b3171501",
         991 => x"13560801",
         992 => x"b356c702",
         993 => x"13150801",
         994 => x"13550501",
         995 => x"3377c702",
         996 => x"b386a602",
         997 => x"93150701",
         998 => x"13d70701",
         999 => x"3367b700",
        1000 => x"637ad700",
        1001 => x"3307e800",
        1002 => x"63660701",
        1003 => x"6374d700",
        1004 => x"33070701",
        1005 => x"3307d740",
        1006 => x"b356c702",
        1007 => x"3377c702",
        1008 => x"b386a602",
        1009 => x"93970701",
        1010 => x"13170701",
        1011 => x"93d70701",
        1012 => x"b3e7e700",
        1013 => x"63fad700",
        1014 => x"b307f800",
        1015 => x"63e60701",
        1016 => x"63f4d700",
        1017 => x"b3870701",
        1018 => x"b387d740",
        1019 => x"33d51701",
        1020 => x"93050000",
        1021 => x"67800000",
        1022 => x"37030001",
        1023 => x"93060001",
        1024 => x"e36666f4",
        1025 => x"93068001",
        1026 => x"6ff05ff4",
        1027 => x"93060000",
        1028 => x"630c0600",
        1029 => x"37070100",
        1030 => x"637ee606",
        1031 => x"93360610",
        1032 => x"93c61600",
        1033 => x"93963600",
        1034 => x"3357d600",
        1035 => x"b388e800",
        1036 => x"03c70800",
        1037 => x"3307d700",
        1038 => x"93060002",
        1039 => x"b388e640",
        1040 => x"6394e606",
        1041 => x"3387c540",
        1042 => x"93550801",
        1043 => x"3356b702",
        1044 => x"13150801",
        1045 => x"13550501",
        1046 => x"93d60701",
        1047 => x"3377b702",
        1048 => x"3306a602",
        1049 => x"13170701",
        1050 => x"33e7e600",
        1051 => x"637ac700",
        1052 => x"3307e800",
        1053 => x"63660701",
        1054 => x"6374c700",
        1055 => x"33070701",
        1056 => x"3307c740",
        1057 => x"b356b702",
        1058 => x"3377b702",
        1059 => x"b386a602",
        1060 => x"6ff05ff3",
        1061 => x"37070001",
        1062 => x"93060001",
        1063 => x"e366e6f8",
        1064 => x"93068001",
        1065 => x"6ff05ff8",
        1066 => x"33181601",
        1067 => x"b3d6e500",
        1068 => x"b3171501",
        1069 => x"b3951501",
        1070 => x"3357e500",
        1071 => x"13550801",
        1072 => x"3367b700",
        1073 => x"b3d5a602",
        1074 => x"13130801",
        1075 => x"13530301",
        1076 => x"b3f6a602",
        1077 => x"b3856502",
        1078 => x"13960601",
        1079 => x"93560701",
        1080 => x"b3e6c600",
        1081 => x"63fab600",
        1082 => x"b306d800",
        1083 => x"63e60601",
        1084 => x"63f4b600",
        1085 => x"b3860601",
        1086 => x"b386b640",
        1087 => x"33d6a602",
        1088 => x"13170701",
        1089 => x"13570701",
        1090 => x"b3f6a602",
        1091 => x"33066602",
        1092 => x"93960601",
        1093 => x"3367d700",
        1094 => x"637ac700",
        1095 => x"3307e800",
        1096 => x"63660701",
        1097 => x"6374c700",
        1098 => x"33070701",
        1099 => x"3307c740",
        1100 => x"6ff09ff1",
        1101 => x"63e4d51c",
        1102 => x"37080100",
        1103 => x"63fe0605",
        1104 => x"13b80610",
        1105 => x"13481800",
        1106 => x"13183800",
        1107 => x"b7380000",
        1108 => x"33d30601",
        1109 => x"938888d3",
        1110 => x"b3886800",
        1111 => x"83c80800",
        1112 => x"13030002",
        1113 => x"b3880801",
        1114 => x"33081341",
        1115 => x"63101305",
        1116 => x"63e4b600",
        1117 => x"636cc500",
        1118 => x"3306c540",
        1119 => x"b386d540",
        1120 => x"3337c500",
        1121 => x"93070600",
        1122 => x"3387e640",
        1123 => x"13850700",
        1124 => x"93050700",
        1125 => x"67800000",
        1126 => x"b7080001",
        1127 => x"13080001",
        1128 => x"e3e616fb",
        1129 => x"13088001",
        1130 => x"6ff05ffa",
        1131 => x"b3571601",
        1132 => x"b3960601",
        1133 => x"b3e6d700",
        1134 => x"33d71501",
        1135 => x"13de0601",
        1136 => x"335fc703",
        1137 => x"13930601",
        1138 => x"13530301",
        1139 => x"b3970501",
        1140 => x"b3551501",
        1141 => x"b3e5f500",
        1142 => x"93d70501",
        1143 => x"33160601",
        1144 => x"33150501",
        1145 => x"3377c703",
        1146 => x"b30ee303",
        1147 => x"13170701",
        1148 => x"b3e7e700",
        1149 => x"13070f00",
        1150 => x"63fed701",
        1151 => x"b387f600",
        1152 => x"1307ffff",
        1153 => x"63e8d700",
        1154 => x"63f6d701",
        1155 => x"1307efff",
        1156 => x"b387d700",
        1157 => x"b387d741",
        1158 => x"b3dec703",
        1159 => x"93950501",
        1160 => x"93d50501",
        1161 => x"b3f7c703",
        1162 => x"138e0e00",
        1163 => x"3303d303",
        1164 => x"93970701",
        1165 => x"b3e5f500",
        1166 => x"63fe6500",
        1167 => x"b385b600",
        1168 => x"138efeff",
        1169 => x"63e8d500",
        1170 => x"63f66500",
        1171 => x"138eeeff",
        1172 => x"b385d500",
        1173 => x"93170701",
        1174 => x"370f0100",
        1175 => x"b3e7c701",
        1176 => x"b3856540",
        1177 => x"1303ffff",
        1178 => x"33f76700",
        1179 => x"135e0601",
        1180 => x"93d70701",
        1181 => x"33736600",
        1182 => x"b30e6702",
        1183 => x"33836702",
        1184 => x"3307c703",
        1185 => x"b387c703",
        1186 => x"330e6700",
        1187 => x"13d70e01",
        1188 => x"3307c701",
        1189 => x"63746700",
        1190 => x"b387e701",
        1191 => x"13530701",
        1192 => x"b307f300",
        1193 => x"37030100",
        1194 => x"1303f3ff",
        1195 => x"33776700",
        1196 => x"13170701",
        1197 => x"b3fe6e00",
        1198 => x"3307d701",
        1199 => x"63e6f500",
        1200 => x"639ef500",
        1201 => x"637ce500",
        1202 => x"3306c740",
        1203 => x"3333c700",
        1204 => x"b306d300",
        1205 => x"13070600",
        1206 => x"b387d740",
        1207 => x"3307e540",
        1208 => x"3335e500",
        1209 => x"b385f540",
        1210 => x"b385a540",
        1211 => x"b3981501",
        1212 => x"33570701",
        1213 => x"33e5e800",
        1214 => x"b3d50501",
        1215 => x"67800000",
        1216 => x"13030500",
        1217 => x"630e0600",
        1218 => x"83830500",
        1219 => x"23007300",
        1220 => x"1306f6ff",
        1221 => x"13031300",
        1222 => x"93851500",
        1223 => x"e31606fe",
        1224 => x"67800000",
        1225 => x"13030500",
        1226 => x"630a0600",
        1227 => x"2300b300",
        1228 => x"1306f6ff",
        1229 => x"13031300",
        1230 => x"e31a06fe",
        1231 => x"67800000",
        1232 => x"630c0602",
        1233 => x"13030500",
        1234 => x"93061000",
        1235 => x"636ab500",
        1236 => x"9306f0ff",
        1237 => x"1307f6ff",
        1238 => x"3303e300",
        1239 => x"b385e500",
        1240 => x"83830500",
        1241 => x"23007300",
        1242 => x"1306f6ff",
        1243 => x"3303d300",
        1244 => x"b385d500",
        1245 => x"e31606fe",
        1246 => x"67800000",
        1247 => x"6f000000",
        1248 => x"130101ff",
        1249 => x"23248100",
        1250 => x"13040000",
        1251 => x"23229100",
        1252 => x"23202101",
        1253 => x"23261100",
        1254 => x"93040500",
        1255 => x"13090400",
        1256 => x"93070400",
        1257 => x"732410c8",
        1258 => x"732910c0",
        1259 => x"f32710c8",
        1260 => x"e31af4fe",
        1261 => x"37460f00",
        1262 => x"13060624",
        1263 => x"93060000",
        1264 => x"13050900",
        1265 => x"93050400",
        1266 => x"eff05fb5",
        1267 => x"37460f00",
        1268 => x"23a4a400",
        1269 => x"93050400",
        1270 => x"13050900",
        1271 => x"13060624",
        1272 => x"93060000",
        1273 => x"eff08ff0",
        1274 => x"8320c100",
        1275 => x"03248100",
        1276 => x"23a0a400",
        1277 => x"23a2b400",
        1278 => x"03290100",
        1279 => x"83244100",
        1280 => x"13050000",
        1281 => x"13010101",
        1282 => x"67800000",
        1283 => x"03a74188",
        1284 => x"b7870020",
        1285 => x"93870700",
        1286 => x"93060040",
        1287 => x"b387d740",
        1288 => x"630c0700",
        1289 => x"3305a700",
        1290 => x"63e2a702",
        1291 => x"23a2a188",
        1292 => x"13050700",
        1293 => x"67800000",
        1294 => x"93868189",
        1295 => x"13878189",
        1296 => x"23a2d188",
        1297 => x"3305a700",
        1298 => x"e3f2a7fe",
        1299 => x"130101ff",
        1300 => x"23261100",
        1301 => x"ef00c03a",
        1302 => x"8320c100",
        1303 => x"9307c000",
        1304 => x"2320f500",
        1305 => x"1307f0ff",
        1306 => x"13050700",
        1307 => x"13010101",
        1308 => x"67800000",
        1309 => x"370700f0",
        1310 => x"83274702",
        1311 => x"93f74700",
        1312 => x"e38c07fe",
        1313 => x"03258702",
        1314 => x"1375f50f",
        1315 => x"67800000",
        1316 => x"b70700f0",
        1317 => x"23a6a702",
        1318 => x"23a0b702",
        1319 => x"67800000",
        1320 => x"1375f50f",
        1321 => x"b70700f0",
        1322 => x"370700f0",
        1323 => x"23a4a702",
        1324 => x"83274702",
        1325 => x"93f70701",
        1326 => x"e38c07fe",
        1327 => x"67800000",
        1328 => x"630e0502",
        1329 => x"130101ff",
        1330 => x"23248100",
        1331 => x"23261100",
        1332 => x"13040500",
        1333 => x"03450500",
        1334 => x"630a0500",
        1335 => x"13041400",
        1336 => x"eff01ffc",
        1337 => x"03450400",
        1338 => x"e31a05fe",
        1339 => x"8320c100",
        1340 => x"03248100",
        1341 => x"13010101",
        1342 => x"67800000",
        1343 => x"67800000",
        1344 => x"130101f9",
        1345 => x"23248106",
        1346 => x"23229106",
        1347 => x"23261106",
        1348 => x"23202107",
        1349 => x"232e3105",
        1350 => x"232c4105",
        1351 => x"232a5105",
        1352 => x"23286105",
        1353 => x"23267105",
        1354 => x"23248105",
        1355 => x"23229105",
        1356 => x"2320a105",
        1357 => x"93040500",
        1358 => x"13840500",
        1359 => x"232c0100",
        1360 => x"232e0100",
        1361 => x"23200102",
        1362 => x"23220102",
        1363 => x"23240102",
        1364 => x"23260102",
        1365 => x"23280102",
        1366 => x"232a0102",
        1367 => x"232c0102",
        1368 => x"232e0102",
        1369 => x"97f2ffff",
        1370 => x"938282d1",
        1371 => x"73905230",
        1372 => x"93050004",
        1373 => x"1305101b",
        1374 => x"eff09ff1",
        1375 => x"37877d01",
        1376 => x"b70700f0",
        1377 => x"1307f783",
        1378 => x"23a6e708",
        1379 => x"93061001",
        1380 => x"37170000",
        1381 => x"23a0d708",
        1382 => x"13077738",
        1383 => x"23a8e70a",
        1384 => x"37270000",
        1385 => x"1307f770",
        1386 => x"23a6e70a",
        1387 => x"23a0d70a",
        1388 => x"13078070",
        1389 => x"23a0e706",
        1390 => x"3707f900",
        1391 => x"13078700",
        1392 => x"23a0e704",
        1393 => x"93020008",
        1394 => x"73904230",
        1395 => x"b7220000",
        1396 => x"93828280",
        1397 => x"73900230",
        1398 => x"b7390000",
        1399 => x"138549e8",
        1400 => x"eff01fee",
        1401 => x"63549002",
        1402 => x"1389f4ff",
        1403 => x"9304f0ff",
        1404 => x"03250400",
        1405 => x"1309f9ff",
        1406 => x"13044400",
        1407 => x"eff05fec",
        1408 => x"138549e8",
        1409 => x"eff0dfeb",
        1410 => x"e31499fe",
        1411 => x"37350000",
        1412 => x"b7faeeee",
        1413 => x"130585e5",
        1414 => x"b7090010",
        1415 => x"37140000",
        1416 => x"1389faee",
        1417 => x"eff0dfe9",
        1418 => x"373b0000",
        1419 => x"9389f9ff",
        1420 => x"938aeaee",
        1421 => x"130404e1",
        1422 => x"93040000",
        1423 => x"b71b0000",
        1424 => x"938b0b2c",
        1425 => x"130af000",
        1426 => x"93050000",
        1427 => x"13058100",
        1428 => x"ef008036",
        1429 => x"938bfbff",
        1430 => x"630a0502",
        1431 => x"e3960bfe",
        1432 => x"73001000",
        1433 => x"b70700f0",
        1434 => x"9306f00f",
        1435 => x"23a4d706",
        1436 => x"03a70704",
        1437 => x"93860704",
        1438 => x"13670730",
        1439 => x"23a0e704",
        1440 => x"93070009",
        1441 => x"23a4f600",
        1442 => x"6ff05ffb",
        1443 => x"032c8100",
        1444 => x"8325c100",
        1445 => x"13060400",
        1446 => x"9357cc01",
        1447 => x"13974500",
        1448 => x"b367f700",
        1449 => x"b3f73701",
        1450 => x"33773c01",
        1451 => x"13d5f541",
        1452 => x"13d88501",
        1453 => x"3307f700",
        1454 => x"33070701",
        1455 => x"9377d500",
        1456 => x"3307f700",
        1457 => x"33774703",
        1458 => x"937725ff",
        1459 => x"93860400",
        1460 => x"13050c00",
        1461 => x"3307f700",
        1462 => x"b307ec40",
        1463 => x"1357f741",
        1464 => x"3338fc00",
        1465 => x"3387e540",
        1466 => x"33070741",
        1467 => x"b3885703",
        1468 => x"33072703",
        1469 => x"33b82703",
        1470 => x"33071701",
        1471 => x"b3872703",
        1472 => x"33070701",
        1473 => x"1358f741",
        1474 => x"13783800",
        1475 => x"b307f800",
        1476 => x"33b80701",
        1477 => x"3307e800",
        1478 => x"1318e701",
        1479 => x"93d72700",
        1480 => x"b367f800",
        1481 => x"13582740",
        1482 => x"93184800",
        1483 => x"13d3c701",
        1484 => x"33e36800",
        1485 => x"33733301",
        1486 => x"b3f83701",
        1487 => x"135e8801",
        1488 => x"1357f741",
        1489 => x"b3886800",
        1490 => x"b388c801",
        1491 => x"1373d700",
        1492 => x"b3886800",
        1493 => x"b3f84803",
        1494 => x"137727ff",
        1495 => x"939c4700",
        1496 => x"b38cfc40",
        1497 => x"939c2c00",
        1498 => x"b30c9c41",
        1499 => x"b388e800",
        1500 => x"33871741",
        1501 => x"93d8f841",
        1502 => x"33b3e700",
        1503 => x"33081841",
        1504 => x"33086840",
        1505 => x"33082803",
        1506 => x"33035703",
        1507 => x"b3382703",
        1508 => x"33086800",
        1509 => x"33072703",
        1510 => x"33081801",
        1511 => x"9358f841",
        1512 => x"93f83800",
        1513 => x"3387e800",
        1514 => x"b3381701",
        1515 => x"b3880801",
        1516 => x"9398e801",
        1517 => x"13572700",
        1518 => x"33e7e800",
        1519 => x"13184700",
        1520 => x"3307e840",
        1521 => x"13172700",
        1522 => x"338de740",
        1523 => x"efe09fea",
        1524 => x"83260101",
        1525 => x"13070500",
        1526 => x"13880c00",
        1527 => x"93070d00",
        1528 => x"13060c00",
        1529 => x"93058be8",
        1530 => x"13058101",
        1531 => x"ef00c015",
        1532 => x"13058101",
        1533 => x"eff0dfcc",
        1534 => x"e3980be4",
        1535 => x"6ff05fe6",
        1536 => x"03a5c187",
        1537 => x"67800000",
        1538 => x"130101ff",
        1539 => x"23248100",
        1540 => x"23261100",
        1541 => x"93070000",
        1542 => x"13040500",
        1543 => x"63880700",
        1544 => x"93050000",
        1545 => x"97000000",
        1546 => x"e7000000",
        1547 => x"b7370000",
        1548 => x"03a587fe",
        1549 => x"83278502",
        1550 => x"63840700",
        1551 => x"e7800700",
        1552 => x"13050400",
        1553 => x"eff09fb3",
        1554 => x"130101ff",
        1555 => x"23248100",
        1556 => x"23229100",
        1557 => x"37340000",
        1558 => x"b7340000",
        1559 => x"9387c4fe",
        1560 => x"1304c4fe",
        1561 => x"3304f440",
        1562 => x"23202101",
        1563 => x"23261100",
        1564 => x"13542440",
        1565 => x"9384c4fe",
        1566 => x"13090000",
        1567 => x"63108904",
        1568 => x"b7340000",
        1569 => x"37340000",
        1570 => x"9387c4fe",
        1571 => x"1304c4fe",
        1572 => x"3304f440",
        1573 => x"13542440",
        1574 => x"9384c4fe",
        1575 => x"13090000",
        1576 => x"63188902",
        1577 => x"8320c100",
        1578 => x"03248100",
        1579 => x"83244100",
        1580 => x"03290100",
        1581 => x"13010101",
        1582 => x"67800000",
        1583 => x"83a70400",
        1584 => x"13091900",
        1585 => x"93844400",
        1586 => x"e7800700",
        1587 => x"6ff01ffb",
        1588 => x"83a70400",
        1589 => x"13091900",
        1590 => x"93844400",
        1591 => x"e7800700",
        1592 => x"6ff01ffc",
        1593 => x"130101f6",
        1594 => x"232af108",
        1595 => x"b7070080",
        1596 => x"93c7f7ff",
        1597 => x"232ef100",
        1598 => x"2328f100",
        1599 => x"b707ffff",
        1600 => x"2326d108",
        1601 => x"2324b100",
        1602 => x"232cb100",
        1603 => x"93878720",
        1604 => x"9306c108",
        1605 => x"93058100",
        1606 => x"232e1106",
        1607 => x"232af100",
        1608 => x"2328e108",
        1609 => x"232c0109",
        1610 => x"232e1109",
        1611 => x"2322d100",
        1612 => x"ef00c040",
        1613 => x"83278100",
        1614 => x"23800700",
        1615 => x"8320c107",
        1616 => x"1301010a",
        1617 => x"67800000",
        1618 => x"130101f6",
        1619 => x"232af108",
        1620 => x"b7070080",
        1621 => x"93c7f7ff",
        1622 => x"232ef100",
        1623 => x"2328f100",
        1624 => x"b707ffff",
        1625 => x"93878720",
        1626 => x"232af100",
        1627 => x"2324a100",
        1628 => x"232ca100",
        1629 => x"03a5c187",
        1630 => x"2324c108",
        1631 => x"2326d108",
        1632 => x"13860500",
        1633 => x"93068108",
        1634 => x"93058100",
        1635 => x"232e1106",
        1636 => x"2328e108",
        1637 => x"232c0109",
        1638 => x"232e1109",
        1639 => x"2322d100",
        1640 => x"ef00c039",
        1641 => x"83278100",
        1642 => x"23800700",
        1643 => x"8320c107",
        1644 => x"1301010a",
        1645 => x"67800000",
        1646 => x"13860500",
        1647 => x"93050500",
        1648 => x"03a5c187",
        1649 => x"6f004000",
        1650 => x"130101ff",
        1651 => x"23248100",
        1652 => x"23229100",
        1653 => x"13040500",
        1654 => x"13850500",
        1655 => x"93050600",
        1656 => x"23261100",
        1657 => x"23a40188",
        1658 => x"eff09f99",
        1659 => x"9307f0ff",
        1660 => x"6318f500",
        1661 => x"83a78188",
        1662 => x"63840700",
        1663 => x"2320f400",
        1664 => x"8320c100",
        1665 => x"03248100",
        1666 => x"83244100",
        1667 => x"13010101",
        1668 => x"67800000",
        1669 => x"130101fe",
        1670 => x"23282101",
        1671 => x"03a98500",
        1672 => x"232c8100",
        1673 => x"23263101",
        1674 => x"23225101",
        1675 => x"23206101",
        1676 => x"232e1100",
        1677 => x"232a9100",
        1678 => x"23244101",
        1679 => x"83aa0500",
        1680 => x"13840500",
        1681 => x"130b0600",
        1682 => x"93890600",
        1683 => x"63ec2609",
        1684 => x"8397c500",
        1685 => x"13f70748",
        1686 => x"63040708",
        1687 => x"03274401",
        1688 => x"93043000",
        1689 => x"83a50501",
        1690 => x"b384e402",
        1691 => x"13072000",
        1692 => x"b38aba40",
        1693 => x"130a0500",
        1694 => x"b3c4e402",
        1695 => x"13871600",
        1696 => x"33075701",
        1697 => x"63f4e400",
        1698 => x"93040700",
        1699 => x"93f70740",
        1700 => x"6386070a",
        1701 => x"93850400",
        1702 => x"13050a00",
        1703 => x"ef001067",
        1704 => x"13090500",
        1705 => x"630c050a",
        1706 => x"83250401",
        1707 => x"13860a00",
        1708 => x"eff01f85",
        1709 => x"8357c400",
        1710 => x"93f7f7b7",
        1711 => x"93e70708",
        1712 => x"2316f400",
        1713 => x"23282401",
        1714 => x"232a9400",
        1715 => x"33095901",
        1716 => x"b3845441",
        1717 => x"23202401",
        1718 => x"23249400",
        1719 => x"13890900",
        1720 => x"63f42901",
        1721 => x"13890900",
        1722 => x"03250400",
        1723 => x"13060900",
        1724 => x"93050b00",
        1725 => x"eff0df84",
        1726 => x"83278400",
        1727 => x"13050000",
        1728 => x"b3872741",
        1729 => x"2324f400",
        1730 => x"83270400",
        1731 => x"b3872701",
        1732 => x"2320f400",
        1733 => x"8320c101",
        1734 => x"03248101",
        1735 => x"83244101",
        1736 => x"03290101",
        1737 => x"8329c100",
        1738 => x"032a8100",
        1739 => x"832a4100",
        1740 => x"032b0100",
        1741 => x"13010102",
        1742 => x"67800000",
        1743 => x"13860400",
        1744 => x"13050a00",
        1745 => x"ef001071",
        1746 => x"13090500",
        1747 => x"e31c05f6",
        1748 => x"83250401",
        1749 => x"13050a00",
        1750 => x"ef00d04b",
        1751 => x"9307c000",
        1752 => x"2320fa00",
        1753 => x"8357c400",
        1754 => x"1305f0ff",
        1755 => x"93e70704",
        1756 => x"2316f400",
        1757 => x"6ff01ffa",
        1758 => x"83278600",
        1759 => x"130101fd",
        1760 => x"232e3101",
        1761 => x"23286101",
        1762 => x"23261102",
        1763 => x"23248102",
        1764 => x"23229102",
        1765 => x"23202103",
        1766 => x"232c4101",
        1767 => x"232a5101",
        1768 => x"23267101",
        1769 => x"23248101",
        1770 => x"23229101",
        1771 => x"2320a101",
        1772 => x"032b0600",
        1773 => x"93090600",
        1774 => x"63940712",
        1775 => x"13050000",
        1776 => x"8320c102",
        1777 => x"03248102",
        1778 => x"23a20900",
        1779 => x"83244102",
        1780 => x"03290102",
        1781 => x"8329c101",
        1782 => x"032a8101",
        1783 => x"832a4101",
        1784 => x"032b0101",
        1785 => x"832bc100",
        1786 => x"032c8100",
        1787 => x"832c4100",
        1788 => x"032d0100",
        1789 => x"13010103",
        1790 => x"67800000",
        1791 => x"832b0b00",
        1792 => x"032d4b00",
        1793 => x"130b8b00",
        1794 => x"03298400",
        1795 => x"832a0400",
        1796 => x"e3060dfe",
        1797 => x"63642d09",
        1798 => x"8317c400",
        1799 => x"13f70748",
        1800 => x"630e0706",
        1801 => x"83244401",
        1802 => x"83250401",
        1803 => x"b3049c02",
        1804 => x"b38aba40",
        1805 => x"13871a00",
        1806 => x"3307a701",
        1807 => x"b3c49403",
        1808 => x"63f4e400",
        1809 => x"93040700",
        1810 => x"93f70740",
        1811 => x"6388070a",
        1812 => x"93850400",
        1813 => x"13050a00",
        1814 => x"ef00504b",
        1815 => x"13090500",
        1816 => x"630e050a",
        1817 => x"83250401",
        1818 => x"13860a00",
        1819 => x"eff04fe9",
        1820 => x"8357c400",
        1821 => x"93f7f7b7",
        1822 => x"93e70708",
        1823 => x"2316f400",
        1824 => x"23282401",
        1825 => x"232a9400",
        1826 => x"33095901",
        1827 => x"b3845441",
        1828 => x"23202401",
        1829 => x"23249400",
        1830 => x"13090d00",
        1831 => x"63742d01",
        1832 => x"13090d00",
        1833 => x"03250400",
        1834 => x"13060900",
        1835 => x"93850b00",
        1836 => x"eff00fe9",
        1837 => x"83278400",
        1838 => x"b3872741",
        1839 => x"2324f400",
        1840 => x"83270400",
        1841 => x"b3872701",
        1842 => x"2320f400",
        1843 => x"83a78900",
        1844 => x"b387a741",
        1845 => x"23a4f900",
        1846 => x"e39207f2",
        1847 => x"6ff01fee",
        1848 => x"130a0500",
        1849 => x"13840500",
        1850 => x"930b0000",
        1851 => x"130d0000",
        1852 => x"130c3000",
        1853 => x"930c2000",
        1854 => x"6ff01ff1",
        1855 => x"13860400",
        1856 => x"13050a00",
        1857 => x"ef001055",
        1858 => x"13090500",
        1859 => x"e31a05f6",
        1860 => x"83250401",
        1861 => x"13050a00",
        1862 => x"ef00d02f",
        1863 => x"9307c000",
        1864 => x"2320fa00",
        1865 => x"8357c400",
        1866 => x"1305f0ff",
        1867 => x"93e70704",
        1868 => x"2316f400",
        1869 => x"23a40900",
        1870 => x"6ff09fe8",
        1871 => x"83d7c500",
        1872 => x"130101f5",
        1873 => x"2324810a",
        1874 => x"2322910a",
        1875 => x"2320210b",
        1876 => x"232c4109",
        1877 => x"2326110a",
        1878 => x"232e3109",
        1879 => x"232a5109",
        1880 => x"23286109",
        1881 => x"23267109",
        1882 => x"23248109",
        1883 => x"23229109",
        1884 => x"2320a109",
        1885 => x"232eb107",
        1886 => x"93f70708",
        1887 => x"130a0500",
        1888 => x"13890500",
        1889 => x"93040600",
        1890 => x"13840600",
        1891 => x"63880706",
        1892 => x"83a70501",
        1893 => x"63940706",
        1894 => x"93050004",
        1895 => x"ef001037",
        1896 => x"2320a900",
        1897 => x"2328a900",
        1898 => x"63160504",
        1899 => x"9307c000",
        1900 => x"2320fa00",
        1901 => x"1305f0ff",
        1902 => x"8320c10a",
        1903 => x"0324810a",
        1904 => x"8324410a",
        1905 => x"0329010a",
        1906 => x"8329c109",
        1907 => x"032a8109",
        1908 => x"832a4109",
        1909 => x"032b0109",
        1910 => x"832bc108",
        1911 => x"032c8108",
        1912 => x"832c4108",
        1913 => x"032d0108",
        1914 => x"832dc107",
        1915 => x"1301010b",
        1916 => x"67800000",
        1917 => x"93070004",
        1918 => x"232af900",
        1919 => x"93070002",
        1920 => x"a304f102",
        1921 => x"93070003",
        1922 => x"23220102",
        1923 => x"2305f102",
        1924 => x"23268100",
        1925 => x"930c5002",
        1926 => x"373b0000",
        1927 => x"b73b0000",
        1928 => x"373d0000",
        1929 => x"372c0000",
        1930 => x"930a0000",
        1931 => x"13840400",
        1932 => x"83470400",
        1933 => x"63840700",
        1934 => x"639c970d",
        1935 => x"b30d9440",
        1936 => x"63069402",
        1937 => x"93860d00",
        1938 => x"13860400",
        1939 => x"93050900",
        1940 => x"13050a00",
        1941 => x"eff01fbc",
        1942 => x"9307f0ff",
        1943 => x"6304f524",
        1944 => x"83274102",
        1945 => x"b387b701",
        1946 => x"2322f102",
        1947 => x"83470400",
        1948 => x"638a0722",
        1949 => x"9307f0ff",
        1950 => x"93041400",
        1951 => x"23280100",
        1952 => x"232e0100",
        1953 => x"232af100",
        1954 => x"232c0100",
        1955 => x"a3090104",
        1956 => x"23240106",
        1957 => x"930d1000",
        1958 => x"83c50400",
        1959 => x"13065000",
        1960 => x"13054bf5",
        1961 => x"ef00d014",
        1962 => x"83270101",
        1963 => x"13841400",
        1964 => x"63140506",
        1965 => x"13f70701",
        1966 => x"63060700",
        1967 => x"13070002",
        1968 => x"a309e104",
        1969 => x"13f78700",
        1970 => x"63060700",
        1971 => x"1307b002",
        1972 => x"a309e104",
        1973 => x"83c60400",
        1974 => x"1307a002",
        1975 => x"638ce604",
        1976 => x"8327c101",
        1977 => x"13840400",
        1978 => x"93060000",
        1979 => x"13069000",
        1980 => x"1305a000",
        1981 => x"03470400",
        1982 => x"93051400",
        1983 => x"130707fd",
        1984 => x"637ee608",
        1985 => x"63840604",
        1986 => x"232ef100",
        1987 => x"6f000004",
        1988 => x"13041400",
        1989 => x"6ff0dff1",
        1990 => x"13074bf5",
        1991 => x"3305e540",
        1992 => x"3395ad00",
        1993 => x"b3e7a700",
        1994 => x"2328f100",
        1995 => x"93040400",
        1996 => x"6ff09ff6",
        1997 => x"0327c100",
        1998 => x"93064700",
        1999 => x"03270700",
        2000 => x"2326d100",
        2001 => x"63420704",
        2002 => x"232ee100",
        2003 => x"03470400",
        2004 => x"9307e002",
        2005 => x"6314f708",
        2006 => x"03471400",
        2007 => x"9307a002",
        2008 => x"6318f704",
        2009 => x"8327c100",
        2010 => x"13042400",
        2011 => x"13874700",
        2012 => x"83a70700",
        2013 => x"2326e100",
        2014 => x"63d40700",
        2015 => x"9307f0ff",
        2016 => x"232af100",
        2017 => x"6f008005",
        2018 => x"3307e040",
        2019 => x"93e72700",
        2020 => x"232ee100",
        2021 => x"2328f100",
        2022 => x"6ff05ffb",
        2023 => x"b387a702",
        2024 => x"13840500",
        2025 => x"93061000",
        2026 => x"b387e700",
        2027 => x"6ff09ff4",
        2028 => x"13041400",
        2029 => x"232a0100",
        2030 => x"93060000",
        2031 => x"93070000",
        2032 => x"13069000",
        2033 => x"1305a000",
        2034 => x"03470400",
        2035 => x"93051400",
        2036 => x"130707fd",
        2037 => x"6372e608",
        2038 => x"e39406fa",
        2039 => x"83450400",
        2040 => x"13063000",
        2041 => x"1385cbf5",
        2042 => x"ef009000",
        2043 => x"63020502",
        2044 => x"9387cbf5",
        2045 => x"3305f540",
        2046 => x"83270101",
        2047 => x"13070004",
        2048 => x"3317a700",
        2049 => x"b3e7e700",
        2050 => x"13041400",
        2051 => x"2328f100",
        2052 => x"83450400",
        2053 => x"13066000",
        2054 => x"13050df6",
        2055 => x"93041400",
        2056 => x"2304b102",
        2057 => x"ef00c07c",
        2058 => x"63080508",
        2059 => x"63980a04",
        2060 => x"03270101",
        2061 => x"8327c100",
        2062 => x"13770710",
        2063 => x"63080702",
        2064 => x"93874700",
        2065 => x"2326f100",
        2066 => x"83274102",
        2067 => x"b3873701",
        2068 => x"2322f102",
        2069 => x"6ff09fdd",
        2070 => x"b387a702",
        2071 => x"13840500",
        2072 => x"93061000",
        2073 => x"b387e700",
        2074 => x"6ff01ff6",
        2075 => x"93877700",
        2076 => x"93f787ff",
        2077 => x"93878700",
        2078 => x"6ff0dffc",
        2079 => x"1307c100",
        2080 => x"93064ca1",
        2081 => x"13060900",
        2082 => x"93050101",
        2083 => x"13050a00",
        2084 => x"97000000",
        2085 => x"e7000000",
        2086 => x"9307f0ff",
        2087 => x"93090500",
        2088 => x"e314f5fa",
        2089 => x"8357c900",
        2090 => x"93f70704",
        2091 => x"e39407d0",
        2092 => x"03254102",
        2093 => x"6ff05fd0",
        2094 => x"1307c100",
        2095 => x"93064ca1",
        2096 => x"13060900",
        2097 => x"93050101",
        2098 => x"13050a00",
        2099 => x"ef00801b",
        2100 => x"6ff09ffc",
        2101 => x"130101fd",
        2102 => x"232a5101",
        2103 => x"83a70501",
        2104 => x"930a0700",
        2105 => x"03a78500",
        2106 => x"23248102",
        2107 => x"23202103",
        2108 => x"232e3101",
        2109 => x"232c4101",
        2110 => x"23261102",
        2111 => x"23229102",
        2112 => x"23286101",
        2113 => x"23267101",
        2114 => x"93090500",
        2115 => x"13840500",
        2116 => x"13090600",
        2117 => x"138a0600",
        2118 => x"63d4e700",
        2119 => x"93070700",
        2120 => x"2320f900",
        2121 => x"03473404",
        2122 => x"63060700",
        2123 => x"93871700",
        2124 => x"2320f900",
        2125 => x"83270400",
        2126 => x"93f70702",
        2127 => x"63880700",
        2128 => x"83270900",
        2129 => x"93872700",
        2130 => x"2320f900",
        2131 => x"83240400",
        2132 => x"93f46400",
        2133 => x"639e0400",
        2134 => x"130b9401",
        2135 => x"930bf0ff",
        2136 => x"8327c400",
        2137 => x"03270900",
        2138 => x"b387e740",
        2139 => x"63c2f408",
        2140 => x"83473404",
        2141 => x"b336f000",
        2142 => x"83270400",
        2143 => x"93f70702",
        2144 => x"6390070c",
        2145 => x"13063404",
        2146 => x"93050a00",
        2147 => x"13850900",
        2148 => x"e7800a00",
        2149 => x"9307f0ff",
        2150 => x"6308f506",
        2151 => x"83270400",
        2152 => x"13074000",
        2153 => x"93040000",
        2154 => x"93f76700",
        2155 => x"639ce700",
        2156 => x"8324c400",
        2157 => x"83270900",
        2158 => x"b384f440",
        2159 => x"63d40400",
        2160 => x"93040000",
        2161 => x"83278400",
        2162 => x"03270401",
        2163 => x"6356f700",
        2164 => x"b387e740",
        2165 => x"b384f400",
        2166 => x"13090000",
        2167 => x"1304a401",
        2168 => x"130bf0ff",
        2169 => x"63902409",
        2170 => x"13050000",
        2171 => x"6f000002",
        2172 => x"93061000",
        2173 => x"13060b00",
        2174 => x"93050a00",
        2175 => x"13850900",
        2176 => x"e7800a00",
        2177 => x"631a7503",
        2178 => x"1305f0ff",
        2179 => x"8320c102",
        2180 => x"03248102",
        2181 => x"83244102",
        2182 => x"03290102",
        2183 => x"8329c101",
        2184 => x"032a8101",
        2185 => x"832a4101",
        2186 => x"032b0101",
        2187 => x"832bc100",
        2188 => x"13010103",
        2189 => x"67800000",
        2190 => x"93841400",
        2191 => x"6ff05ff2",
        2192 => x"3307d400",
        2193 => x"13060003",
        2194 => x"a301c704",
        2195 => x"03475404",
        2196 => x"93871600",
        2197 => x"b307f400",
        2198 => x"93862600",
        2199 => x"a381e704",
        2200 => x"6ff05ff2",
        2201 => x"93061000",
        2202 => x"13060400",
        2203 => x"93050a00",
        2204 => x"13850900",
        2205 => x"e7800a00",
        2206 => x"e30865f9",
        2207 => x"13091900",
        2208 => x"6ff05ff6",
        2209 => x"130101fd",
        2210 => x"23248102",
        2211 => x"23229102",
        2212 => x"23202103",
        2213 => x"232e3101",
        2214 => x"23261102",
        2215 => x"232c4101",
        2216 => x"232a5101",
        2217 => x"23286101",
        2218 => x"83c88501",
        2219 => x"93078007",
        2220 => x"93040500",
        2221 => x"13840500",
        2222 => x"13090600",
        2223 => x"93890600",
        2224 => x"63ee1701",
        2225 => x"93072006",
        2226 => x"93863504",
        2227 => x"63ee1701",
        2228 => x"638a082a",
        2229 => x"93078005",
        2230 => x"638af820",
        2231 => x"930a2404",
        2232 => x"23011405",
        2233 => x"6f004004",
        2234 => x"9387d8f9",
        2235 => x"93f7f70f",
        2236 => x"13065001",
        2237 => x"e364f6fe",
        2238 => x"37360000",
        2239 => x"93972700",
        2240 => x"130606f9",
        2241 => x"b387c700",
        2242 => x"83a70700",
        2243 => x"67800700",
        2244 => x"83270700",
        2245 => x"938a2504",
        2246 => x"93864700",
        2247 => x"83a70700",
        2248 => x"2320d700",
        2249 => x"2381f504",
        2250 => x"93071000",
        2251 => x"6f004029",
        2252 => x"03a60500",
        2253 => x"83270700",
        2254 => x"13750608",
        2255 => x"93854700",
        2256 => x"630e0504",
        2257 => x"83a70700",
        2258 => x"2320b700",
        2259 => x"37370000",
        2260 => x"83254400",
        2261 => x"130887f6",
        2262 => x"63d2071e",
        2263 => x"1307d002",
        2264 => x"a301e404",
        2265 => x"2324b400",
        2266 => x"63d80504",
        2267 => x"b307f040",
        2268 => x"1307a000",
        2269 => x"938a0600",
        2270 => x"33f6e702",
        2271 => x"938afaff",
        2272 => x"3306c800",
        2273 => x"03460600",
        2274 => x"2380ca00",
        2275 => x"13860700",
        2276 => x"b3d7e702",
        2277 => x"e372e6fe",
        2278 => x"6f008009",
        2279 => x"83a70700",
        2280 => x"13750604",
        2281 => x"2320b700",
        2282 => x"e30205fa",
        2283 => x"93970701",
        2284 => x"93d70741",
        2285 => x"6ff09ff9",
        2286 => x"1376b6ff",
        2287 => x"2320c400",
        2288 => x"6ff0dffa",
        2289 => x"03a60500",
        2290 => x"83270700",
        2291 => x"13750608",
        2292 => x"93854700",
        2293 => x"63080500",
        2294 => x"2320b700",
        2295 => x"83a70700",
        2296 => x"6f004001",
        2297 => x"13760604",
        2298 => x"2320b700",
        2299 => x"e30806fe",
        2300 => x"83d70700",
        2301 => x"37380000",
        2302 => x"1307f006",
        2303 => x"130888f6",
        2304 => x"639ae812",
        2305 => x"13078000",
        2306 => x"a3010404",
        2307 => x"03264400",
        2308 => x"2324c400",
        2309 => x"e34006f6",
        2310 => x"83250400",
        2311 => x"93f5b5ff",
        2312 => x"2320b400",
        2313 => x"e39807f4",
        2314 => x"938a0600",
        2315 => x"e31406f4",
        2316 => x"93078000",
        2317 => x"6314f702",
        2318 => x"83270400",
        2319 => x"93f71700",
        2320 => x"638e0700",
        2321 => x"03274400",
        2322 => x"83270401",
        2323 => x"63c8e700",
        2324 => x"93070003",
        2325 => x"a38ffafe",
        2326 => x"938afaff",
        2327 => x"b3865641",
        2328 => x"2328d400",
        2329 => x"13870900",
        2330 => x"93060900",
        2331 => x"1306c100",
        2332 => x"93050400",
        2333 => x"13850400",
        2334 => x"eff0dfc5",
        2335 => x"130af0ff",
        2336 => x"63164515",
        2337 => x"1305f0ff",
        2338 => x"8320c102",
        2339 => x"03248102",
        2340 => x"83244102",
        2341 => x"03290102",
        2342 => x"8329c101",
        2343 => x"032a8101",
        2344 => x"832a4101",
        2345 => x"032b0101",
        2346 => x"13010103",
        2347 => x"67800000",
        2348 => x"83a70500",
        2349 => x"93e70702",
        2350 => x"23a0f500",
        2351 => x"37380000",
        2352 => x"93088007",
        2353 => x"1308c8f7",
        2354 => x"03260400",
        2355 => x"a3021405",
        2356 => x"83270700",
        2357 => x"13750608",
        2358 => x"93854700",
        2359 => x"630e0500",
        2360 => x"2320b700",
        2361 => x"83a70700",
        2362 => x"6f000002",
        2363 => x"37380000",
        2364 => x"130888f6",
        2365 => x"6ff05ffd",
        2366 => x"13750604",
        2367 => x"2320b700",
        2368 => x"e30205fe",
        2369 => x"83d70700",
        2370 => x"13771600",
        2371 => x"63060700",
        2372 => x"13660602",
        2373 => x"2320c400",
        2374 => x"63860700",
        2375 => x"13070001",
        2376 => x"6ff09fee",
        2377 => x"03270400",
        2378 => x"1377f7fd",
        2379 => x"2320e400",
        2380 => x"6ff0dffe",
        2381 => x"1307a000",
        2382 => x"6ff01fed",
        2383 => x"130887f6",
        2384 => x"1307a000",
        2385 => x"6ff09fec",
        2386 => x"03a60500",
        2387 => x"83270700",
        2388 => x"83a54501",
        2389 => x"13780608",
        2390 => x"13854700",
        2391 => x"630a0800",
        2392 => x"2320a700",
        2393 => x"83a70700",
        2394 => x"23a0b700",
        2395 => x"6f008001",
        2396 => x"2320a700",
        2397 => x"13760604",
        2398 => x"83a70700",
        2399 => x"e30606fe",
        2400 => x"2390b700",
        2401 => x"23280400",
        2402 => x"938a0600",
        2403 => x"6ff09fed",
        2404 => x"83270700",
        2405 => x"03a64500",
        2406 => x"93050000",
        2407 => x"93864700",
        2408 => x"2320d700",
        2409 => x"83aa0700",
        2410 => x"13850a00",
        2411 => x"ef004024",
        2412 => x"63060500",
        2413 => x"33055541",
        2414 => x"2322a400",
        2415 => x"83274400",
        2416 => x"2328f400",
        2417 => x"a3010404",
        2418 => x"6ff0dfe9",
        2419 => x"83260401",
        2420 => x"13860a00",
        2421 => x"93050900",
        2422 => x"13850400",
        2423 => x"e7800900",
        2424 => x"e30245eb",
        2425 => x"83270400",
        2426 => x"93f72700",
        2427 => x"63940704",
        2428 => x"8327c100",
        2429 => x"0325c400",
        2430 => x"e358f5e8",
        2431 => x"13850700",
        2432 => x"6ff09fe8",
        2433 => x"93061000",
        2434 => x"13860a00",
        2435 => x"93050900",
        2436 => x"13850400",
        2437 => x"e7800900",
        2438 => x"e30665e7",
        2439 => x"130a1a00",
        2440 => x"8327c400",
        2441 => x"0327c100",
        2442 => x"b387e740",
        2443 => x"e34cfafc",
        2444 => x"6ff01ffc",
        2445 => x"130a0000",
        2446 => x"930a9401",
        2447 => x"130bf0ff",
        2448 => x"6ff01ffe",
        2449 => x"130101ff",
        2450 => x"23248100",
        2451 => x"13840500",
        2452 => x"83a50500",
        2453 => x"23229100",
        2454 => x"23261100",
        2455 => x"93040500",
        2456 => x"63840500",
        2457 => x"eff01ffe",
        2458 => x"93050400",
        2459 => x"03248100",
        2460 => x"8320c100",
        2461 => x"13850400",
        2462 => x"83244100",
        2463 => x"13010101",
        2464 => x"6f004019",
        2465 => x"83a7c187",
        2466 => x"6382a716",
        2467 => x"83274502",
        2468 => x"130101fe",
        2469 => x"232c8100",
        2470 => x"232e1100",
        2471 => x"232a9100",
        2472 => x"23282101",
        2473 => x"23263101",
        2474 => x"13040500",
        2475 => x"638a0704",
        2476 => x"83a7c700",
        2477 => x"638c0702",
        2478 => x"93040000",
        2479 => x"13090008",
        2480 => x"83274402",
        2481 => x"83a7c700",
        2482 => x"b3879700",
        2483 => x"83a50700",
        2484 => x"6396050e",
        2485 => x"93844400",
        2486 => x"e39424ff",
        2487 => x"83274402",
        2488 => x"13050400",
        2489 => x"83a5c700",
        2490 => x"ef00c012",
        2491 => x"83274402",
        2492 => x"83a50700",
        2493 => x"63860500",
        2494 => x"13050400",
        2495 => x"ef008011",
        2496 => x"83254401",
        2497 => x"63860500",
        2498 => x"13050400",
        2499 => x"ef008010",
        2500 => x"83254402",
        2501 => x"63860500",
        2502 => x"13050400",
        2503 => x"ef00800f",
        2504 => x"83258403",
        2505 => x"63860500",
        2506 => x"13050400",
        2507 => x"ef00800e",
        2508 => x"8325c403",
        2509 => x"63860500",
        2510 => x"13050400",
        2511 => x"ef00800d",
        2512 => x"83250404",
        2513 => x"63860500",
        2514 => x"13050400",
        2515 => x"ef00800c",
        2516 => x"8325c405",
        2517 => x"63860500",
        2518 => x"13050400",
        2519 => x"ef00800b",
        2520 => x"83258405",
        2521 => x"63860500",
        2522 => x"13050400",
        2523 => x"ef00800a",
        2524 => x"83254403",
        2525 => x"63860500",
        2526 => x"13050400",
        2527 => x"ef008009",
        2528 => x"83278401",
        2529 => x"63860704",
        2530 => x"83278402",
        2531 => x"13050400",
        2532 => x"e7800700",
        2533 => x"83258404",
        2534 => x"638c0502",
        2535 => x"13050400",
        2536 => x"03248101",
        2537 => x"8320c101",
        2538 => x"83244101",
        2539 => x"03290101",
        2540 => x"8329c100",
        2541 => x"13010102",
        2542 => x"6ff0dfe8",
        2543 => x"83a90500",
        2544 => x"13050400",
        2545 => x"ef000005",
        2546 => x"93850900",
        2547 => x"6ff05ff0",
        2548 => x"8320c101",
        2549 => x"03248101",
        2550 => x"83244101",
        2551 => x"03290101",
        2552 => x"8329c100",
        2553 => x"13010102",
        2554 => x"67800000",
        2555 => x"67800000",
        2556 => x"93f5f50f",
        2557 => x"3306c500",
        2558 => x"6316c500",
        2559 => x"13050000",
        2560 => x"67800000",
        2561 => x"83470500",
        2562 => x"e38cb7fe",
        2563 => x"13051500",
        2564 => x"6ff09ffe",
        2565 => x"638a050e",
        2566 => x"83a7c5ff",
        2567 => x"130101fe",
        2568 => x"232c8100",
        2569 => x"232e1100",
        2570 => x"1384c5ff",
        2571 => x"63d40700",
        2572 => x"3304f400",
        2573 => x"2326a100",
        2574 => x"ef008033",
        2575 => x"83a70189",
        2576 => x"0325c100",
        2577 => x"639e0700",
        2578 => x"23220400",
        2579 => x"23a88188",
        2580 => x"03248101",
        2581 => x"8320c101",
        2582 => x"13010102",
        2583 => x"6f008031",
        2584 => x"6374f402",
        2585 => x"03260400",
        2586 => x"b306c400",
        2587 => x"639ad700",
        2588 => x"83a60700",
        2589 => x"83a74700",
        2590 => x"b386c600",
        2591 => x"2320d400",
        2592 => x"2322f400",
        2593 => x"6ff09ffc",
        2594 => x"13870700",
        2595 => x"83a74700",
        2596 => x"63840700",
        2597 => x"e37af4fe",
        2598 => x"83260700",
        2599 => x"3306d700",
        2600 => x"63188602",
        2601 => x"03260400",
        2602 => x"b386c600",
        2603 => x"2320d700",
        2604 => x"3306d700",
        2605 => x"e39ec7f8",
        2606 => x"03a60700",
        2607 => x"83a74700",
        2608 => x"b306d600",
        2609 => x"2320d700",
        2610 => x"2322f700",
        2611 => x"6ff05ff8",
        2612 => x"6378c400",
        2613 => x"9307c000",
        2614 => x"2320f500",
        2615 => x"6ff05ff7",
        2616 => x"03260400",
        2617 => x"b306c400",
        2618 => x"639ad700",
        2619 => x"83a60700",
        2620 => x"83a74700",
        2621 => x"b386c600",
        2622 => x"2320d400",
        2623 => x"2322f400",
        2624 => x"23228700",
        2625 => x"6ff0dff4",
        2626 => x"67800000",
        2627 => x"130101fe",
        2628 => x"232a9100",
        2629 => x"93843500",
        2630 => x"93f4c4ff",
        2631 => x"23282101",
        2632 => x"232e1100",
        2633 => x"232c8100",
        2634 => x"23263101",
        2635 => x"93848400",
        2636 => x"9307c000",
        2637 => x"13090500",
        2638 => x"63f0f406",
        2639 => x"9304c000",
        2640 => x"63eeb404",
        2641 => x"13050900",
        2642 => x"ef008022",
        2643 => x"03a70189",
        2644 => x"13040700",
        2645 => x"63180406",
        2646 => x"83a7c188",
        2647 => x"639a0700",
        2648 => x"93050000",
        2649 => x"13050900",
        2650 => x"ef00001c",
        2651 => x"23a6a188",
        2652 => x"93850400",
        2653 => x"13050900",
        2654 => x"ef00001b",
        2655 => x"9309f0ff",
        2656 => x"631a350b",
        2657 => x"9307c000",
        2658 => x"2320f900",
        2659 => x"13050900",
        2660 => x"ef00401e",
        2661 => x"6f000001",
        2662 => x"e3d404fa",
        2663 => x"9307c000",
        2664 => x"2320f900",
        2665 => x"13050000",
        2666 => x"8320c101",
        2667 => x"03248101",
        2668 => x"83244101",
        2669 => x"03290101",
        2670 => x"8329c100",
        2671 => x"13010102",
        2672 => x"67800000",
        2673 => x"83270400",
        2674 => x"b3879740",
        2675 => x"63ce0704",
        2676 => x"1306b000",
        2677 => x"637af600",
        2678 => x"2320f400",
        2679 => x"3304f400",
        2680 => x"23209400",
        2681 => x"6f000001",
        2682 => x"83274400",
        2683 => x"631a8702",
        2684 => x"23a8f188",
        2685 => x"13050900",
        2686 => x"ef00c017",
        2687 => x"1305b400",
        2688 => x"93074400",
        2689 => x"137585ff",
        2690 => x"3307f540",
        2691 => x"e30ef5f8",
        2692 => x"3304e400",
        2693 => x"b387a740",
        2694 => x"2320f400",
        2695 => x"6ff0dff8",
        2696 => x"2322f700",
        2697 => x"6ff01ffd",
        2698 => x"13070400",
        2699 => x"03244400",
        2700 => x"6ff05ff2",
        2701 => x"13043500",
        2702 => x"1374c4ff",
        2703 => x"e30285fa",
        2704 => x"b305a440",
        2705 => x"13050900",
        2706 => x"ef00000e",
        2707 => x"e31a35f9",
        2708 => x"6ff05ff3",
        2709 => x"130101fe",
        2710 => x"232c8100",
        2711 => x"232e1100",
        2712 => x"232a9100",
        2713 => x"23282101",
        2714 => x"23263101",
        2715 => x"23244101",
        2716 => x"13040600",
        2717 => x"63940502",
        2718 => x"03248101",
        2719 => x"8320c101",
        2720 => x"83244101",
        2721 => x"03290101",
        2722 => x"8329c100",
        2723 => x"032a8100",
        2724 => x"93050600",
        2725 => x"13010102",
        2726 => x"6ff05fe7",
        2727 => x"63180602",
        2728 => x"eff05fd7",
        2729 => x"93040000",
        2730 => x"8320c101",
        2731 => x"03248101",
        2732 => x"03290101",
        2733 => x"8329c100",
        2734 => x"032a8100",
        2735 => x"13850400",
        2736 => x"83244101",
        2737 => x"13010102",
        2738 => x"67800000",
        2739 => x"130a0500",
        2740 => x"93840500",
        2741 => x"ef00400a",
        2742 => x"13090500",
        2743 => x"63668500",
        2744 => x"93571500",
        2745 => x"e3e287fc",
        2746 => x"93050400",
        2747 => x"13050a00",
        2748 => x"eff0dfe1",
        2749 => x"93090500",
        2750 => x"e30605fa",
        2751 => x"13060400",
        2752 => x"63748900",
        2753 => x"13060900",
        2754 => x"93850400",
        2755 => x"13850900",
        2756 => x"efe00fff",
        2757 => x"93850400",
        2758 => x"13050a00",
        2759 => x"eff09fcf",
        2760 => x"93840900",
        2761 => x"6ff05ff8",
        2762 => x"130101ff",
        2763 => x"23248100",
        2764 => x"23229100",
        2765 => x"13040500",
        2766 => x"13850500",
        2767 => x"23261100",
        2768 => x"23a40188",
        2769 => x"efe09f8c",
        2770 => x"9307f0ff",
        2771 => x"6318f500",
        2772 => x"83a78188",
        2773 => x"63840700",
        2774 => x"2320f400",
        2775 => x"8320c100",
        2776 => x"03248100",
        2777 => x"83244100",
        2778 => x"13010101",
        2779 => x"67800000",
        2780 => x"67800000",
        2781 => x"67800000",
        2782 => x"83a7c5ff",
        2783 => x"1385c7ff",
        2784 => x"63d80700",
        2785 => x"b385a500",
        2786 => x"83a70500",
        2787 => x"3305f500",
        2788 => x"67800000",
        2789 => x"10000000",
        2790 => x"00000000",
        2791 => x"037a5200",
        2792 => x"017c0101",
        2793 => x"1b0d0200",
        2794 => x"10000000",
        2795 => x"18000000",
        2796 => x"c4daffff",
        2797 => x"78040000",
        2798 => x"00000000",
        2799 => x"10000000",
        2800 => x"00000000",
        2801 => x"037a5200",
        2802 => x"017c0101",
        2803 => x"1b0d0200",
        2804 => x"10000000",
        2805 => x"18000000",
        2806 => x"14dfffff",
        2807 => x"30040000",
        2808 => x"00000000",
        2809 => x"10000000",
        2810 => x"00000000",
        2811 => x"037a5200",
        2812 => x"017c0101",
        2813 => x"1b0d0200",
        2814 => x"10000000",
        2815 => x"18000000",
        2816 => x"1ce3ffff",
        2817 => x"e4030000",
        2818 => x"00000000",
        2819 => x"30313233",
        2820 => x"34353637",
        2821 => x"38396162",
        2822 => x"63646566",
        2823 => x"00000000",
        2824 => x"58040000",
        2825 => x"64040000",
        2826 => x"34040000",
        2827 => x"4c040000",
        2828 => x"40040000",
        2829 => x"74030000",
        2830 => x"74030000",
        2831 => x"74030000",
        2832 => x"a8040000",
        2833 => x"74030000",
        2834 => x"74030000",
        2835 => x"74030000",
        2836 => x"74030000",
        2837 => x"74030000",
        2838 => x"74030000",
        2839 => x"74030000",
        2840 => x"70040000",
        2841 => x"0c050000",
        2842 => x"c4040000",
        2843 => x"c4040000",
        2844 => x"c4040000",
        2845 => x"c4040000",
        2846 => x"00050000",
        2847 => x"4c050000",
        2848 => x"24050000",
        2849 => x"c4040000",
        2850 => x"c4040000",
        2851 => x"c4040000",
        2852 => x"c4040000",
        2853 => x"c4040000",
        2854 => x"c4040000",
        2855 => x"c4040000",
        2856 => x"c4040000",
        2857 => x"c4040000",
        2858 => x"c4040000",
        2859 => x"c4040000",
        2860 => x"c4040000",
        2861 => x"c4040000",
        2862 => x"c4040000",
        2863 => x"ec040000",
        2864 => x"ec040000",
        2865 => x"c4040000",
        2866 => x"c4040000",
        2867 => x"c4040000",
        2868 => x"c4040000",
        2869 => x"c4040000",
        2870 => x"c4040000",
        2871 => x"c4040000",
        2872 => x"c4040000",
        2873 => x"c4040000",
        2874 => x"c4040000",
        2875 => x"c4040000",
        2876 => x"c4040000",
        2877 => x"00050000",
        2878 => x"0c050000",
        2879 => x"c8050000",
        2880 => x"b0050000",
        2881 => x"c4040000",
        2882 => x"c4040000",
        2883 => x"c4040000",
        2884 => x"c4040000",
        2885 => x"c4040000",
        2886 => x"c4040000",
        2887 => x"98050000",
        2888 => x"c4040000",
        2889 => x"c4040000",
        2890 => x"c4040000",
        2891 => x"c4040000",
        2892 => x"ec040000",
        2893 => x"ec040000",
        2894 => x"00010202",
        2895 => x"03030303",
        2896 => x"04040404",
        2897 => x"04040404",
        2898 => x"05050505",
        2899 => x"05050505",
        2900 => x"05050505",
        2901 => x"05050505",
        2902 => x"06060606",
        2903 => x"06060606",
        2904 => x"06060606",
        2905 => x"06060606",
        2906 => x"06060606",
        2907 => x"06060606",
        2908 => x"06060606",
        2909 => x"06060606",
        2910 => x"07070707",
        2911 => x"07070707",
        2912 => x"07070707",
        2913 => x"07070707",
        2914 => x"07070707",
        2915 => x"07070707",
        2916 => x"07070707",
        2917 => x"07070707",
        2918 => x"07070707",
        2919 => x"07070707",
        2920 => x"07070707",
        2921 => x"07070707",
        2922 => x"07070707",
        2923 => x"07070707",
        2924 => x"07070707",
        2925 => x"07070707",
        2926 => x"08080808",
        2927 => x"08080808",
        2928 => x"08080808",
        2929 => x"08080808",
        2930 => x"08080808",
        2931 => x"08080808",
        2932 => x"08080808",
        2933 => x"08080808",
        2934 => x"08080808",
        2935 => x"08080808",
        2936 => x"08080808",
        2937 => x"08080808",
        2938 => x"08080808",
        2939 => x"08080808",
        2940 => x"08080808",
        2941 => x"08080808",
        2942 => x"08080808",
        2943 => x"08080808",
        2944 => x"08080808",
        2945 => x"08080808",
        2946 => x"08080808",
        2947 => x"08080808",
        2948 => x"08080808",
        2949 => x"08080808",
        2950 => x"08080808",
        2951 => x"08080808",
        2952 => x"08080808",
        2953 => x"08080808",
        2954 => x"08080808",
        2955 => x"08080808",
        2956 => x"08080808",
        2957 => x"08080808",
        2958 => x"0d0a4542",
        2959 => x"5245414b",
        2960 => x"21206d65",
        2961 => x"7063203d",
        2962 => x"20000000",
        2963 => x"20696e73",
        2964 => x"6e203d20",
        2965 => x"00000000",
        2966 => x"0d0a0d0a",
        2967 => x"44697370",
        2968 => x"6c617969",
        2969 => x"6e672074",
        2970 => x"68652074",
        2971 => x"696d6520",
        2972 => x"70617373",
        2973 => x"65642073",
        2974 => x"696e6365",
        2975 => x"20726573",
        2976 => x"65740d0a",
        2977 => x"0d0a0000",
        2978 => x"2530356c",
        2979 => x"643a2530",
        2980 => x"366c6420",
        2981 => x"20202530",
        2982 => x"326c643a",
        2983 => x"2530326c",
        2984 => x"643a2530",
        2985 => x"326c640d",
        2986 => x"00000000",
        2987 => x"696e7465",
        2988 => x"72727570",
        2989 => x"745f6469",
        2990 => x"72656374",
        2991 => x"00000000",
        2992 => x"54485541",
        2993 => x"53205249",
        2994 => x"53432d56",
        2995 => x"20525633",
        2996 => x"32494d20",
        2997 => x"62617265",
        2998 => x"206d6574",
        2999 => x"616c2070",
        3000 => x"726f6365",
        3001 => x"73736f72",
        3002 => x"00000000",
        3003 => x"54686520",
        3004 => x"48616775",
        3005 => x"6520556e",
        3006 => x"69766572",
        3007 => x"73697479",
        3008 => x"206f6620",
        3009 => x"4170706c",
        3010 => x"69656420",
        3011 => x"53636965",
        3012 => x"6e636573",
        3013 => x"00000000",
        3014 => x"44657061",
        3015 => x"72746d65",
        3016 => x"6e74206f",
        3017 => x"6620456c",
        3018 => x"65637472",
        3019 => x"6963616c",
        3020 => x"20456e67",
        3021 => x"696e6565",
        3022 => x"72696e67",
        3023 => x"00000000",
        3024 => x"4a2e452e",
        3025 => x"4a2e206f",
        3026 => x"70206465",
        3027 => x"6e204272",
        3028 => x"6f757700",
        3029 => x"232d302b",
        3030 => x"20000000",
        3031 => x"686c4c00",
        3032 => x"65666745",
        3033 => x"46470000",
        3034 => x"30313233",
        3035 => x"34353637",
        3036 => x"38394142",
        3037 => x"43444546",
        3038 => x"00000000",
        3039 => x"30313233",
        3040 => x"34353637",
        3041 => x"38396162",
        3042 => x"63646566",
        3043 => x"00000000",
        3044 => x"10230000",
        3045 => x"30230000",
        3046 => x"dc220000",
        3047 => x"dc220000",
        3048 => x"dc220000",
        3049 => x"dc220000",
        3050 => x"30230000",
        3051 => x"dc220000",
        3052 => x"dc220000",
        3053 => x"dc220000",
        3054 => x"dc220000",
        3055 => x"48250000",
        3056 => x"c4230000",
        3057 => x"b0240000",
        3058 => x"dc220000",
        3059 => x"dc220000",
        3060 => x"90250000",
        3061 => x"dc220000",
        3062 => x"c4230000",
        3063 => x"dc220000",
        3064 => x"dc220000",
        3065 => x"bc240000",
        3066 => x"18000020",
        3067 => x"ac2e0000",
        3068 => x"c02e0000",
        3069 => x"ec2e0000",
        3070 => x"182f0000",
        3071 => x"402f0000",
        3072 => x"00000000",
        3073 => x"00000000",
        3074 => x"00000000",
        3075 => x"00000000",
        3076 => x"00000000",
        3077 => x"00000000",
        3078 => x"00000000",
        3079 => x"00000000",
        3080 => x"00000000",
        3081 => x"00000000",
        3082 => x"00000000",
        3083 => x"00000000",
        3084 => x"00000000",
        3085 => x"00000000",
        3086 => x"00000000",
        3087 => x"00000000",
        3088 => x"00000000",
        3089 => x"00000000",
        3090 => x"00000000",
        3091 => x"00000000",
        3092 => x"00000000",
        3093 => x"00000000",
        3094 => x"00000000",
        3095 => x"00000000",
        3096 => x"00000000",
        3097 => x"80000020",
        3098 => x"18000020",
        others => (others => '0')
    );
end package processor_common_rom;
