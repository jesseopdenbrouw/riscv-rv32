-- srec2vhdl table generator
-- for input file interrupt_direct.srec

library ieee;
use ieee.std_logic_1164.all;

library work;
use work.processor_common.all;

package processor_common_rom is
    constant rom_contents : rom_type := (
           0 => x"97020000",
           1 => x"93828226",
           2 => x"73905230",
           3 => x"97010020",
           4 => x"9381417f",
           5 => x"17810020",
           6 => x"1301c1fe",
           7 => x"13860188",
           8 => x"93874189",
           9 => x"637af600",
          10 => x"3386c740",
          11 => x"93050000",
          12 => x"13850188",
          13 => x"ef10c035",
          14 => x"37050020",
          15 => x"13060500",
          16 => x"93870188",
          17 => x"637cf600",
          18 => x"b7350000",
          19 => x"3386c740",
          20 => x"938585fc",
          21 => x"13050500",
          22 => x"ef104031",
          23 => x"ef10c07c",
          24 => x"b7050020",
          25 => x"13060000",
          26 => x"93850500",
          27 => x"13055000",
          28 => x"ef100047",
          29 => x"ef104077",
          30 => x"6f00c05d",
          31 => x"130101ff",
          32 => x"23261100",
          33 => x"ef00c05f",
          34 => x"8320c100",
          35 => x"13051000",
          36 => x"13010101",
          37 => x"67800000",
          38 => x"130101fd",
          39 => x"232c4101",
          40 => x"130a0500",
          41 => x"37350000",
          42 => x"130545e1",
          43 => x"23248102",
          44 => x"23229102",
          45 => x"23202103",
          46 => x"232e3101",
          47 => x"83244a08",
          48 => x"23261102",
          49 => x"13044100",
          50 => x"ef00805d",
          51 => x"37390000",
          52 => x"9309c1ff",
          53 => x"93070400",
          54 => x"1309c9be",
          55 => x"13f7f400",
          56 => x"3307e900",
          57 => x"03470700",
          58 => x"9387f7ff",
          59 => x"93d44400",
          60 => x"2384e700",
          61 => x"e39437ff",
          62 => x"13054100",
          63 => x"23060100",
          64 => x"ef00005a",
          65 => x"37350000",
          66 => x"130585e2",
          67 => x"ef004059",
          68 => x"03278a08",
          69 => x"9377f700",
          70 => x"b307f900",
          71 => x"83c70700",
          72 => x"1304f4ff",
          73 => x"13574700",
          74 => x"2304f400",
          75 => x"e31434ff",
          76 => x"13054100",
          77 => x"ef00c056",
          78 => x"37350000",
          79 => x"130505e6",
          80 => x"ef000056",
          81 => x"8320c102",
          82 => x"03248102",
          83 => x"83244102",
          84 => x"03290102",
          85 => x"8329c101",
          86 => x"032a8101",
          87 => x"13010103",
          88 => x"67800000",
          89 => x"b70700f0",
          90 => x"03a74708",
          91 => x"1377f7fe",
          92 => x"23a2e708",
          93 => x"03a74700",
          94 => x"13471700",
          95 => x"23a2e700",
          96 => x"67800000",
          97 => x"370700f0",
          98 => x"83274700",
          99 => x"93e70720",
         100 => x"2322f700",
         101 => x"6f000000",
         102 => x"b70700f0",
         103 => x"83a6470f",
         104 => x"03a6070f",
         105 => x"03a7470f",
         106 => x"e31ad7fe",
         107 => x"b7860100",
         108 => x"9305f0ff",
         109 => x"9386066a",
         110 => x"23aeb70e",
         111 => x"b306d600",
         112 => x"23acb70e",
         113 => x"33b6c600",
         114 => x"23acd70e",
         115 => x"3306e600",
         116 => x"23aec70e",
         117 => x"03a74700",
         118 => x"13472700",
         119 => x"23a2e700",
         120 => x"67800000",
         121 => x"b70700f0",
         122 => x"03a74702",
         123 => x"13774700",
         124 => x"630a0700",
         125 => x"03a74700",
         126 => x"13478700",
         127 => x"23a2e700",
         128 => x"83a78702",
         129 => x"67800000",
         130 => x"b70700f0",
         131 => x"03a7470a",
         132 => x"1377f7f0",
         133 => x"23a2e70a",
         134 => x"03a74700",
         135 => x"13474700",
         136 => x"23a2e700",
         137 => x"67800000",
         138 => x"b70700f0",
         139 => x"03a74706",
         140 => x"137777ff",
         141 => x"23a2e706",
         142 => x"03a74700",
         143 => x"13470701",
         144 => x"23a2e700",
         145 => x"67800000",
         146 => x"b70700f0",
         147 => x"03a74704",
         148 => x"137777fe",
         149 => x"23a2e704",
         150 => x"03a74700",
         151 => x"13470702",
         152 => x"23a2e700",
         153 => x"67800000",
         154 => x"6f000000",
         155 => x"13050000",
         156 => x"67800000",
         157 => x"13050000",
         158 => x"67800000",
         159 => x"130101f7",
         160 => x"23221100",
         161 => x"23242100",
         162 => x"23263100",
         163 => x"23284100",
         164 => x"232a5100",
         165 => x"232c6100",
         166 => x"232e7100",
         167 => x"23208102",
         168 => x"23229102",
         169 => x"2324a102",
         170 => x"2326b102",
         171 => x"2328c102",
         172 => x"232ad102",
         173 => x"232ce102",
         174 => x"232ef102",
         175 => x"23200105",
         176 => x"23221105",
         177 => x"23242105",
         178 => x"23263105",
         179 => x"23284105",
         180 => x"232a5105",
         181 => x"232c6105",
         182 => x"232e7105",
         183 => x"23208107",
         184 => x"23229107",
         185 => x"2324a107",
         186 => x"2326b107",
         187 => x"2328c107",
         188 => x"232ad107",
         189 => x"232ce107",
         190 => x"232ef107",
         191 => x"f3222034",
         192 => x"23205108",
         193 => x"f3221034",
         194 => x"23225108",
         195 => x"83a20200",
         196 => x"23245108",
         197 => x"f3223034",
         198 => x"23265108",
         199 => x"f3272034",
         200 => x"37070080",
         201 => x"93067700",
         202 => x"6386d70e",
         203 => x"9306b000",
         204 => x"63fef602",
         205 => x"9346f7fe",
         206 => x"b386d700",
         207 => x"13064000",
         208 => x"636ad602",
         209 => x"1347e7fe",
         210 => x"b387e700",
         211 => x"13073000",
         212 => x"6364f714",
         213 => x"37370000",
         214 => x"93972700",
         215 => x"130707c0",
         216 => x"b387e700",
         217 => x"83a70700",
         218 => x"67800700",
         219 => x"13071000",
         220 => x"6364f708",
         221 => x"03258102",
         222 => x"832fc107",
         223 => x"032f8107",
         224 => x"832e4107",
         225 => x"032e0107",
         226 => x"832dc106",
         227 => x"032d8106",
         228 => x"832c4106",
         229 => x"032c0106",
         230 => x"832bc105",
         231 => x"032b8105",
         232 => x"832a4105",
         233 => x"032a0105",
         234 => x"8329c104",
         235 => x"03298104",
         236 => x"83284104",
         237 => x"03280104",
         238 => x"8327c103",
         239 => x"03278103",
         240 => x"83264103",
         241 => x"03260103",
         242 => x"8325c102",
         243 => x"83244102",
         244 => x"03240102",
         245 => x"8323c101",
         246 => x"03238101",
         247 => x"83224101",
         248 => x"03220101",
         249 => x"8321c100",
         250 => x"03218100",
         251 => x"83204100",
         252 => x"13010109",
         253 => x"73002030",
         254 => x"e3eef6f6",
         255 => x"37370000",
         256 => x"93972700",
         257 => x"130707c1",
         258 => x"b387e700",
         259 => x"83a70700",
         260 => x"67800700",
         261 => x"eff05fd8",
         262 => x"03258102",
         263 => x"6ff0dff5",
         264 => x"eff09fde",
         265 => x"03258102",
         266 => x"6ff01ff5",
         267 => x"eff0dfdf",
         268 => x"03258102",
         269 => x"6ff05ff4",
         270 => x"eff01fe1",
         271 => x"03258102",
         272 => x"6ff09ff3",
         273 => x"eff01fda",
         274 => x"03258102",
         275 => x"6ff0dff2",
         276 => x"9307600d",
         277 => x"6384f806",
         278 => x"9307900a",
         279 => x"6388f818",
         280 => x"63ca170f",
         281 => x"938878fc",
         282 => x"93074002",
         283 => x"63ec1703",
         284 => x"b7370000",
         285 => x"938707c4",
         286 => x"93982800",
         287 => x"b388f800",
         288 => x"83a70800",
         289 => x"67800700",
         290 => x"13050100",
         291 => x"eff0dfc0",
         292 => x"03258102",
         293 => x"6ff05fee",
         294 => x"eff0dfcc",
         295 => x"03258102",
         296 => x"6ff09fed",
         297 => x"ef10c033",
         298 => x"93078005",
         299 => x"2320f500",
         300 => x"9307f0ff",
         301 => x"13850700",
         302 => x"6ff01fec",
         303 => x"63120510",
         304 => x"13858189",
         305 => x"13050500",
         306 => x"6ff01feb",
         307 => x"b7270000",
         308 => x"23a2f500",
         309 => x"93070000",
         310 => x"13850700",
         311 => x"6ff0dfe9",
         312 => x"93070000",
         313 => x"13850700",
         314 => x"6ff01fe9",
         315 => x"ef10402f",
         316 => x"93079000",
         317 => x"2320f500",
         318 => x"9307f0ff",
         319 => x"13850700",
         320 => x"6ff09fe7",
         321 => x"13090600",
         322 => x"13840500",
         323 => x"635cc000",
         324 => x"b384c500",
         325 => x"03450400",
         326 => x"13041400",
         327 => x"eff01fb6",
         328 => x"e39a84fe",
         329 => x"13050900",
         330 => x"6ff01fe5",
         331 => x"13090600",
         332 => x"13840500",
         333 => x"e358c0fe",
         334 => x"b384c500",
         335 => x"eff0dfb3",
         336 => x"2300a400",
         337 => x"13041400",
         338 => x"e31a94fe",
         339 => x"13050900",
         340 => x"6ff09fe2",
         341 => x"938808c0",
         342 => x"9307f000",
         343 => x"e3e417f5",
         344 => x"b7370000",
         345 => x"938747cd",
         346 => x"93982800",
         347 => x"b388f800",
         348 => x"83a70800",
         349 => x"67800700",
         350 => x"ef108026",
         351 => x"9307d000",
         352 => x"2320f500",
         353 => x"9307f0ff",
         354 => x"13850700",
         355 => x"6ff0dfde",
         356 => x"ef100025",
         357 => x"93072000",
         358 => x"2320f500",
         359 => x"9307f0ff",
         360 => x"13850700",
         361 => x"6ff05fdd",
         362 => x"ef108023",
         363 => x"9307f001",
         364 => x"2320f500",
         365 => x"9307f0ff",
         366 => x"13850700",
         367 => x"6ff0dfdb",
         368 => x"b7870020",
         369 => x"93870700",
         370 => x"13070040",
         371 => x"b387e740",
         372 => x"e36af5ee",
         373 => x"ef10c020",
         374 => x"9307c000",
         375 => x"2320f500",
         376 => x"1305f0ff",
         377 => x"13050500",
         378 => x"6ff01fd9",
         379 => x"13090000",
         380 => x"93040500",
         381 => x"13040900",
         382 => x"93090900",
         383 => x"93070900",
         384 => x"732410c8",
         385 => x"f32910c0",
         386 => x"f32710c8",
         387 => x"e31af4fe",
         388 => x"37460f00",
         389 => x"13060624",
         390 => x"93060000",
         391 => x"13850900",
         392 => x"93050400",
         393 => x"ef005016",
         394 => x"37460f00",
         395 => x"23a4a400",
         396 => x"13060624",
         397 => x"93060000",
         398 => x"13850900",
         399 => x"93050400",
         400 => x"ef008051",
         401 => x"23a0a400",
         402 => x"23a2b400",
         403 => x"13050900",
         404 => x"6ff09fd2",
         405 => x"370700f0",
         406 => x"83274702",
         407 => x"93f74700",
         408 => x"e38c07fe",
         409 => x"03258702",
         410 => x"1375f50f",
         411 => x"67800000",
         412 => x"b70700f0",
         413 => x"23a6a702",
         414 => x"23a0b702",
         415 => x"67800000",
         416 => x"1375f50f",
         417 => x"b70700f0",
         418 => x"370700f0",
         419 => x"23a4a702",
         420 => x"83274702",
         421 => x"93f70701",
         422 => x"e38c07fe",
         423 => x"67800000",
         424 => x"630e0502",
         425 => x"130101ff",
         426 => x"23248100",
         427 => x"23261100",
         428 => x"13040500",
         429 => x"03450500",
         430 => x"630a0500",
         431 => x"13041400",
         432 => x"eff01ffc",
         433 => x"03450400",
         434 => x"e31a05fe",
         435 => x"8320c100",
         436 => x"03248100",
         437 => x"13010101",
         438 => x"67800000",
         439 => x"67800000",
         440 => x"13030500",
         441 => x"138e0500",
         442 => x"93080000",
         443 => x"63dc0500",
         444 => x"b337a000",
         445 => x"330eb040",
         446 => x"330efe40",
         447 => x"3303a040",
         448 => x"9308f0ff",
         449 => x"63dc0600",
         450 => x"b337c000",
         451 => x"b306d040",
         452 => x"93c8f8ff",
         453 => x"b386f640",
         454 => x"3306c040",
         455 => x"13070600",
         456 => x"13080300",
         457 => x"93070e00",
         458 => x"639c0628",
         459 => x"b7350000",
         460 => x"938545d1",
         461 => x"6376ce0e",
         462 => x"b7060100",
         463 => x"6378d60c",
         464 => x"93360610",
         465 => x"93c61600",
         466 => x"93963600",
         467 => x"3355d600",
         468 => x"b385a500",
         469 => x"83c50500",
         470 => x"13050002",
         471 => x"b386d500",
         472 => x"b305d540",
         473 => x"630cd500",
         474 => x"b317be00",
         475 => x"b356d300",
         476 => x"3317b600",
         477 => x"b3e7f600",
         478 => x"3318b300",
         479 => x"93550701",
         480 => x"33deb702",
         481 => x"13160701",
         482 => x"13560601",
         483 => x"b3f7b702",
         484 => x"13050e00",
         485 => x"3303c603",
         486 => x"93960701",
         487 => x"93570801",
         488 => x"b3e7d700",
         489 => x"63fe6700",
         490 => x"b307f700",
         491 => x"1305feff",
         492 => x"63e8e700",
         493 => x"63f66700",
         494 => x"1305eeff",
         495 => x"b387e700",
         496 => x"b3876740",
         497 => x"33d3b702",
         498 => x"13180801",
         499 => x"13580801",
         500 => x"b3f7b702",
         501 => x"b3066602",
         502 => x"93970701",
         503 => x"3368f800",
         504 => x"93070300",
         505 => x"637cd800",
         506 => x"33080701",
         507 => x"9307f3ff",
         508 => x"6366e800",
         509 => x"6374d800",
         510 => x"9307e3ff",
         511 => x"13150501",
         512 => x"3365f500",
         513 => x"93050000",
         514 => x"6f00000e",
         515 => x"37050001",
         516 => x"93060001",
         517 => x"e36ca6f2",
         518 => x"93068001",
         519 => x"6ff01ff3",
         520 => x"93060000",
         521 => x"630c0600",
         522 => x"b7070100",
         523 => x"637af60c",
         524 => x"93360610",
         525 => x"93c61600",
         526 => x"93963600",
         527 => x"b357d600",
         528 => x"b385f500",
         529 => x"83c70500",
         530 => x"b387d700",
         531 => x"93060002",
         532 => x"b385f640",
         533 => x"6390f60c",
         534 => x"b307ce40",
         535 => x"93051000",
         536 => x"13530701",
         537 => x"b3de6702",
         538 => x"13160701",
         539 => x"13560601",
         540 => x"93560801",
         541 => x"b3f76702",
         542 => x"13850e00",
         543 => x"330ed603",
         544 => x"93970701",
         545 => x"b3e7f600",
         546 => x"63fec701",
         547 => x"b307f700",
         548 => x"1385feff",
         549 => x"63e8e700",
         550 => x"63f6c701",
         551 => x"1385eeff",
         552 => x"b387e700",
         553 => x"b387c741",
         554 => x"33de6702",
         555 => x"13180801",
         556 => x"13580801",
         557 => x"b3f76702",
         558 => x"b306c603",
         559 => x"93970701",
         560 => x"3368f800",
         561 => x"93070e00",
         562 => x"637cd800",
         563 => x"33080701",
         564 => x"9307feff",
         565 => x"6366e800",
         566 => x"6374d800",
         567 => x"9307eeff",
         568 => x"13150501",
         569 => x"3365f500",
         570 => x"638a0800",
         571 => x"b337a000",
         572 => x"b305b040",
         573 => x"b385f540",
         574 => x"3305a040",
         575 => x"67800000",
         576 => x"b7070001",
         577 => x"93060001",
         578 => x"e36af6f2",
         579 => x"93068001",
         580 => x"6ff0dff2",
         581 => x"3317b600",
         582 => x"b356fe00",
         583 => x"13550701",
         584 => x"331ebe00",
         585 => x"b357f300",
         586 => x"b3e7c701",
         587 => x"33dea602",
         588 => x"13160701",
         589 => x"13560601",
         590 => x"3318b300",
         591 => x"b3f6a602",
         592 => x"3303c603",
         593 => x"93950601",
         594 => x"93d60701",
         595 => x"b3e6b600",
         596 => x"93050e00",
         597 => x"63fe6600",
         598 => x"b306d700",
         599 => x"9305feff",
         600 => x"63e8e600",
         601 => x"63f66600",
         602 => x"9305eeff",
         603 => x"b386e600",
         604 => x"b3866640",
         605 => x"33d3a602",
         606 => x"93970701",
         607 => x"93d70701",
         608 => x"b3f6a602",
         609 => x"33066602",
         610 => x"93960601",
         611 => x"b3e7d700",
         612 => x"93060300",
         613 => x"63fec700",
         614 => x"b307f700",
         615 => x"9306f3ff",
         616 => x"63e8e700",
         617 => x"63f6c700",
         618 => x"9306e3ff",
         619 => x"b387e700",
         620 => x"93950501",
         621 => x"b387c740",
         622 => x"b3e5d500",
         623 => x"6ff05fea",
         624 => x"6366de18",
         625 => x"b7070100",
         626 => x"63f4f604",
         627 => x"13b70610",
         628 => x"13471700",
         629 => x"13173700",
         630 => x"b7370000",
         631 => x"b3d5e600",
         632 => x"938747d1",
         633 => x"b387b700",
         634 => x"83c70700",
         635 => x"b387e700",
         636 => x"13070002",
         637 => x"b305f740",
         638 => x"6316f702",
         639 => x"13051000",
         640 => x"e3e4c6ef",
         641 => x"3335c300",
         642 => x"13451500",
         643 => x"6ff0dfed",
         644 => x"b7070001",
         645 => x"13070001",
         646 => x"e3e0f6fc",
         647 => x"13078001",
         648 => x"6ff09ffb",
         649 => x"3357f600",
         650 => x"b396b600",
         651 => x"b366d700",
         652 => x"3357fe00",
         653 => x"331ebe00",
         654 => x"b357f300",
         655 => x"b3e7c701",
         656 => x"13de0601",
         657 => x"335fc703",
         658 => x"13980601",
         659 => x"13580801",
         660 => x"3316b600",
         661 => x"3377c703",
         662 => x"b30ee803",
         663 => x"13150701",
         664 => x"13d70701",
         665 => x"3367a700",
         666 => x"13050f00",
         667 => x"637ed701",
         668 => x"3387e600",
         669 => x"1305ffff",
         670 => x"6368d700",
         671 => x"6376d701",
         672 => x"1305efff",
         673 => x"3307d700",
         674 => x"3307d741",
         675 => x"b35ec703",
         676 => x"93970701",
         677 => x"93d70701",
         678 => x"3377c703",
         679 => x"3308d803",
         680 => x"13170701",
         681 => x"b3e7e700",
         682 => x"13870e00",
         683 => x"63fe0701",
         684 => x"b387f600",
         685 => x"1387feff",
         686 => x"63e8d700",
         687 => x"63f60701",
         688 => x"1387eeff",
         689 => x"b387d700",
         690 => x"13150501",
         691 => x"b70e0100",
         692 => x"3365e500",
         693 => x"9386feff",
         694 => x"3377d500",
         695 => x"b3870741",
         696 => x"b376d600",
         697 => x"13580501",
         698 => x"13560601",
         699 => x"330ed702",
         700 => x"b306d802",
         701 => x"3307c702",
         702 => x"3308c802",
         703 => x"3306d700",
         704 => x"13570e01",
         705 => x"3307c700",
         706 => x"6374d700",
         707 => x"3308d801",
         708 => x"93560701",
         709 => x"b3860601",
         710 => x"63e6d702",
         711 => x"e394d7ce",
         712 => x"b7070100",
         713 => x"9387f7ff",
         714 => x"3377f700",
         715 => x"13170701",
         716 => x"337efe00",
         717 => x"3313b300",
         718 => x"3307c701",
         719 => x"93050000",
         720 => x"e374e3da",
         721 => x"1305f5ff",
         722 => x"6ff0dfcb",
         723 => x"93050000",
         724 => x"13050000",
         725 => x"6ff05fd9",
         726 => x"93080500",
         727 => x"13830500",
         728 => x"13070600",
         729 => x"13080500",
         730 => x"93870500",
         731 => x"63920628",
         732 => x"b7350000",
         733 => x"938545d1",
         734 => x"6376c30e",
         735 => x"b7060100",
         736 => x"6378d60c",
         737 => x"93360610",
         738 => x"93c61600",
         739 => x"93963600",
         740 => x"3355d600",
         741 => x"b385a500",
         742 => x"83c50500",
         743 => x"13050002",
         744 => x"b386d500",
         745 => x"b305d540",
         746 => x"630cd500",
         747 => x"b317b300",
         748 => x"b3d6d800",
         749 => x"3317b600",
         750 => x"b3e7f600",
         751 => x"3398b800",
         752 => x"93550701",
         753 => x"33d3b702",
         754 => x"13160701",
         755 => x"13560601",
         756 => x"b3f7b702",
         757 => x"13050300",
         758 => x"b3086602",
         759 => x"93960701",
         760 => x"93570801",
         761 => x"b3e7d700",
         762 => x"63fe1701",
         763 => x"b307f700",
         764 => x"1305f3ff",
         765 => x"63e8e700",
         766 => x"63f61701",
         767 => x"1305e3ff",
         768 => x"b387e700",
         769 => x"b3871741",
         770 => x"b3d8b702",
         771 => x"13180801",
         772 => x"13580801",
         773 => x"b3f7b702",
         774 => x"b3061603",
         775 => x"93970701",
         776 => x"3368f800",
         777 => x"93870800",
         778 => x"637cd800",
         779 => x"33080701",
         780 => x"9387f8ff",
         781 => x"6366e800",
         782 => x"6374d800",
         783 => x"9387e8ff",
         784 => x"13150501",
         785 => x"3365f500",
         786 => x"93050000",
         787 => x"67800000",
         788 => x"37050001",
         789 => x"93060001",
         790 => x"e36ca6f2",
         791 => x"93068001",
         792 => x"6ff01ff3",
         793 => x"93060000",
         794 => x"630c0600",
         795 => x"b7070100",
         796 => x"6370f60c",
         797 => x"93360610",
         798 => x"93c61600",
         799 => x"93963600",
         800 => x"b357d600",
         801 => x"b385f500",
         802 => x"83c70500",
         803 => x"b387d700",
         804 => x"93060002",
         805 => x"b385f640",
         806 => x"6396f60a",
         807 => x"b307c340",
         808 => x"93051000",
         809 => x"93580701",
         810 => x"33de1703",
         811 => x"13160701",
         812 => x"13560601",
         813 => x"93560801",
         814 => x"b3f71703",
         815 => x"13050e00",
         816 => x"3303c603",
         817 => x"93970701",
         818 => x"b3e7f600",
         819 => x"63fe6700",
         820 => x"b307f700",
         821 => x"1305feff",
         822 => x"63e8e700",
         823 => x"63f66700",
         824 => x"1305eeff",
         825 => x"b387e700",
         826 => x"b3876740",
         827 => x"33d31703",
         828 => x"13180801",
         829 => x"13580801",
         830 => x"b3f71703",
         831 => x"b3066602",
         832 => x"93970701",
         833 => x"3368f800",
         834 => x"93070300",
         835 => x"637cd800",
         836 => x"33080701",
         837 => x"9307f3ff",
         838 => x"6366e800",
         839 => x"6374d800",
         840 => x"9307e3ff",
         841 => x"13150501",
         842 => x"3365f500",
         843 => x"67800000",
         844 => x"b7070001",
         845 => x"93060001",
         846 => x"e364f6f4",
         847 => x"93068001",
         848 => x"6ff01ff4",
         849 => x"3317b600",
         850 => x"b356f300",
         851 => x"13550701",
         852 => x"3313b300",
         853 => x"b3d7f800",
         854 => x"b3e76700",
         855 => x"33d3a602",
         856 => x"13160701",
         857 => x"13560601",
         858 => x"3398b800",
         859 => x"b3f6a602",
         860 => x"b3086602",
         861 => x"93950601",
         862 => x"93d60701",
         863 => x"b3e6b600",
         864 => x"93050300",
         865 => x"63fe1601",
         866 => x"b306d700",
         867 => x"9305f3ff",
         868 => x"63e8e600",
         869 => x"63f61601",
         870 => x"9305e3ff",
         871 => x"b386e600",
         872 => x"b3861641",
         873 => x"b3d8a602",
         874 => x"93970701",
         875 => x"93d70701",
         876 => x"b3f6a602",
         877 => x"33061603",
         878 => x"93960601",
         879 => x"b3e7d700",
         880 => x"93860800",
         881 => x"63fec700",
         882 => x"b307f700",
         883 => x"9386f8ff",
         884 => x"63e8e700",
         885 => x"63f6c700",
         886 => x"9386e8ff",
         887 => x"b387e700",
         888 => x"93950501",
         889 => x"b387c740",
         890 => x"b3e5d500",
         891 => x"6ff09feb",
         892 => x"63e6d518",
         893 => x"b7070100",
         894 => x"63f4f604",
         895 => x"13b70610",
         896 => x"13471700",
         897 => x"13173700",
         898 => x"b7370000",
         899 => x"b3d5e600",
         900 => x"938747d1",
         901 => x"b387b700",
         902 => x"83c70700",
         903 => x"b387e700",
         904 => x"13070002",
         905 => x"b305f740",
         906 => x"6316f702",
         907 => x"13051000",
         908 => x"e3ee66e0",
         909 => x"33b5c800",
         910 => x"13451500",
         911 => x"67800000",
         912 => x"b7070001",
         913 => x"13070001",
         914 => x"e3e0f6fc",
         915 => x"13078001",
         916 => x"6ff09ffb",
         917 => x"3357f600",
         918 => x"b396b600",
         919 => x"b366d700",
         920 => x"3357f300",
         921 => x"3313b300",
         922 => x"b3d7f800",
         923 => x"b3e76700",
         924 => x"13d30601",
         925 => x"b35e6702",
         926 => x"13980601",
         927 => x"13580801",
         928 => x"3316b600",
         929 => x"33776702",
         930 => x"330ed803",
         931 => x"13150701",
         932 => x"13d70701",
         933 => x"3367a700",
         934 => x"13850e00",
         935 => x"637ec701",
         936 => x"3387e600",
         937 => x"1385feff",
         938 => x"6368d700",
         939 => x"6376c701",
         940 => x"1385eeff",
         941 => x"3307d700",
         942 => x"3307c741",
         943 => x"335e6702",
         944 => x"93970701",
         945 => x"93d70701",
         946 => x"33776702",
         947 => x"3308c803",
         948 => x"13170701",
         949 => x"b3e7e700",
         950 => x"13070e00",
         951 => x"63fe0701",
         952 => x"b387f600",
         953 => x"1307feff",
         954 => x"63e8d700",
         955 => x"63f60701",
         956 => x"1307eeff",
         957 => x"b387d700",
         958 => x"13150501",
         959 => x"370e0100",
         960 => x"3365e500",
         961 => x"9306feff",
         962 => x"3377d500",
         963 => x"b3870741",
         964 => x"b376d600",
         965 => x"13580501",
         966 => x"13560601",
         967 => x"3303d702",
         968 => x"b306d802",
         969 => x"3307c702",
         970 => x"3308c802",
         971 => x"3306d700",
         972 => x"13570301",
         973 => x"3307c700",
         974 => x"6374d700",
         975 => x"3308c801",
         976 => x"93560701",
         977 => x"b3860601",
         978 => x"63e6d702",
         979 => x"e39ed7ce",
         980 => x"b7070100",
         981 => x"9387f7ff",
         982 => x"3377f700",
         983 => x"13170701",
         984 => x"3373f300",
         985 => x"b398b800",
         986 => x"33076700",
         987 => x"93050000",
         988 => x"e3fee8cc",
         989 => x"1305f5ff",
         990 => x"6ff01fcd",
         991 => x"93050000",
         992 => x"13050000",
         993 => x"67800000",
         994 => x"13080600",
         995 => x"93070500",
         996 => x"13870500",
         997 => x"63960620",
         998 => x"b7380000",
         999 => x"938848d1",
        1000 => x"63fcc50c",
        1001 => x"b7060100",
        1002 => x"637ed60a",
        1003 => x"93360610",
        1004 => x"93c61600",
        1005 => x"93963600",
        1006 => x"3353d600",
        1007 => x"b3886800",
        1008 => x"83c80800",
        1009 => x"13030002",
        1010 => x"b386d800",
        1011 => x"b308d340",
        1012 => x"630cd300",
        1013 => x"33971501",
        1014 => x"b356d500",
        1015 => x"33181601",
        1016 => x"33e7e600",
        1017 => x"b3171501",
        1018 => x"13560801",
        1019 => x"b356c702",
        1020 => x"13150801",
        1021 => x"13550501",
        1022 => x"3377c702",
        1023 => x"b386a602",
        1024 => x"93150701",
        1025 => x"13d70701",
        1026 => x"3367b700",
        1027 => x"637ad700",
        1028 => x"3307e800",
        1029 => x"63660701",
        1030 => x"6374d700",
        1031 => x"33070701",
        1032 => x"3307d740",
        1033 => x"b356c702",
        1034 => x"3377c702",
        1035 => x"b386a602",
        1036 => x"93970701",
        1037 => x"13170701",
        1038 => x"93d70701",
        1039 => x"b3e7e700",
        1040 => x"63fad700",
        1041 => x"b307f800",
        1042 => x"63e60701",
        1043 => x"63f4d700",
        1044 => x"b3870701",
        1045 => x"b387d740",
        1046 => x"33d51701",
        1047 => x"93050000",
        1048 => x"67800000",
        1049 => x"37030001",
        1050 => x"93060001",
        1051 => x"e36666f4",
        1052 => x"93068001",
        1053 => x"6ff05ff4",
        1054 => x"93060000",
        1055 => x"630c0600",
        1056 => x"37070100",
        1057 => x"637ee606",
        1058 => x"93360610",
        1059 => x"93c61600",
        1060 => x"93963600",
        1061 => x"3357d600",
        1062 => x"b388e800",
        1063 => x"03c70800",
        1064 => x"3307d700",
        1065 => x"93060002",
        1066 => x"b388e640",
        1067 => x"6394e606",
        1068 => x"3387c540",
        1069 => x"93550801",
        1070 => x"3356b702",
        1071 => x"13150801",
        1072 => x"13550501",
        1073 => x"93d60701",
        1074 => x"3377b702",
        1075 => x"3306a602",
        1076 => x"13170701",
        1077 => x"33e7e600",
        1078 => x"637ac700",
        1079 => x"3307e800",
        1080 => x"63660701",
        1081 => x"6374c700",
        1082 => x"33070701",
        1083 => x"3307c740",
        1084 => x"b356b702",
        1085 => x"3377b702",
        1086 => x"b386a602",
        1087 => x"6ff05ff3",
        1088 => x"37070001",
        1089 => x"93060001",
        1090 => x"e366e6f8",
        1091 => x"93068001",
        1092 => x"6ff05ff8",
        1093 => x"33181601",
        1094 => x"b3d6e500",
        1095 => x"b3171501",
        1096 => x"b3951501",
        1097 => x"3357e500",
        1098 => x"13550801",
        1099 => x"3367b700",
        1100 => x"b3d5a602",
        1101 => x"13130801",
        1102 => x"13530301",
        1103 => x"b3f6a602",
        1104 => x"b3856502",
        1105 => x"13960601",
        1106 => x"93560701",
        1107 => x"b3e6c600",
        1108 => x"63fab600",
        1109 => x"b306d800",
        1110 => x"63e60601",
        1111 => x"63f4b600",
        1112 => x"b3860601",
        1113 => x"b386b640",
        1114 => x"33d6a602",
        1115 => x"13170701",
        1116 => x"13570701",
        1117 => x"b3f6a602",
        1118 => x"33066602",
        1119 => x"93960601",
        1120 => x"3367d700",
        1121 => x"637ac700",
        1122 => x"3307e800",
        1123 => x"63660701",
        1124 => x"6374c700",
        1125 => x"33070701",
        1126 => x"3307c740",
        1127 => x"6ff09ff1",
        1128 => x"63e4d51c",
        1129 => x"37080100",
        1130 => x"63fe0605",
        1131 => x"13b80610",
        1132 => x"13481800",
        1133 => x"13183800",
        1134 => x"b7380000",
        1135 => x"33d30601",
        1136 => x"938848d1",
        1137 => x"b3886800",
        1138 => x"83c80800",
        1139 => x"13030002",
        1140 => x"b3880801",
        1141 => x"33081341",
        1142 => x"63101305",
        1143 => x"63e4b600",
        1144 => x"636cc500",
        1145 => x"3306c540",
        1146 => x"b386d540",
        1147 => x"3337c500",
        1148 => x"93070600",
        1149 => x"3387e640",
        1150 => x"13850700",
        1151 => x"93050700",
        1152 => x"67800000",
        1153 => x"b7080001",
        1154 => x"13080001",
        1155 => x"e3e616fb",
        1156 => x"13088001",
        1157 => x"6ff05ffa",
        1158 => x"b3571601",
        1159 => x"b3960601",
        1160 => x"b3e6d700",
        1161 => x"33d71501",
        1162 => x"13de0601",
        1163 => x"335fc703",
        1164 => x"13930601",
        1165 => x"13530301",
        1166 => x"b3970501",
        1167 => x"b3551501",
        1168 => x"b3e5f500",
        1169 => x"93d70501",
        1170 => x"33160601",
        1171 => x"33150501",
        1172 => x"3377c703",
        1173 => x"b30ee303",
        1174 => x"13170701",
        1175 => x"b3e7e700",
        1176 => x"13070f00",
        1177 => x"63fed701",
        1178 => x"b387f600",
        1179 => x"1307ffff",
        1180 => x"63e8d700",
        1181 => x"63f6d701",
        1182 => x"1307efff",
        1183 => x"b387d700",
        1184 => x"b387d741",
        1185 => x"b3dec703",
        1186 => x"93950501",
        1187 => x"93d50501",
        1188 => x"b3f7c703",
        1189 => x"138e0e00",
        1190 => x"3303d303",
        1191 => x"93970701",
        1192 => x"b3e5f500",
        1193 => x"63fe6500",
        1194 => x"b385b600",
        1195 => x"138efeff",
        1196 => x"63e8d500",
        1197 => x"63f66500",
        1198 => x"138eeeff",
        1199 => x"b385d500",
        1200 => x"93170701",
        1201 => x"370f0100",
        1202 => x"b3e7c701",
        1203 => x"b3856540",
        1204 => x"1303ffff",
        1205 => x"33f76700",
        1206 => x"135e0601",
        1207 => x"93d70701",
        1208 => x"33736600",
        1209 => x"b30e6702",
        1210 => x"33836702",
        1211 => x"3307c703",
        1212 => x"b387c703",
        1213 => x"330e6700",
        1214 => x"13d70e01",
        1215 => x"3307c701",
        1216 => x"63746700",
        1217 => x"b387e701",
        1218 => x"13530701",
        1219 => x"b307f300",
        1220 => x"37030100",
        1221 => x"1303f3ff",
        1222 => x"33776700",
        1223 => x"13170701",
        1224 => x"b3fe6e00",
        1225 => x"3307d701",
        1226 => x"63e6f500",
        1227 => x"639ef500",
        1228 => x"637ce500",
        1229 => x"3306c740",
        1230 => x"3333c700",
        1231 => x"b306d300",
        1232 => x"13070600",
        1233 => x"b387d740",
        1234 => x"3307e540",
        1235 => x"3335e500",
        1236 => x"b385f540",
        1237 => x"b385a540",
        1238 => x"b3981501",
        1239 => x"33570701",
        1240 => x"33e5e800",
        1241 => x"b3d50501",
        1242 => x"67800000",
        1243 => x"13030500",
        1244 => x"630e0600",
        1245 => x"83830500",
        1246 => x"23007300",
        1247 => x"1306f6ff",
        1248 => x"13031300",
        1249 => x"93851500",
        1250 => x"e31606fe",
        1251 => x"67800000",
        1252 => x"13030500",
        1253 => x"630a0600",
        1254 => x"2300b300",
        1255 => x"1306f6ff",
        1256 => x"13031300",
        1257 => x"e31a06fe",
        1258 => x"67800000",
        1259 => x"630c0602",
        1260 => x"13030500",
        1261 => x"93061000",
        1262 => x"636ab500",
        1263 => x"9306f0ff",
        1264 => x"1307f6ff",
        1265 => x"3303e300",
        1266 => x"b385e500",
        1267 => x"83830500",
        1268 => x"23007300",
        1269 => x"1306f6ff",
        1270 => x"3303d300",
        1271 => x"b385d500",
        1272 => x"e31606fe",
        1273 => x"67800000",
        1274 => x"6f000000",
        1275 => x"130101ff",
        1276 => x"23248100",
        1277 => x"13040000",
        1278 => x"23229100",
        1279 => x"23202101",
        1280 => x"23261100",
        1281 => x"93040500",
        1282 => x"13090400",
        1283 => x"93070400",
        1284 => x"732410c8",
        1285 => x"732910c0",
        1286 => x"f32710c8",
        1287 => x"e31af4fe",
        1288 => x"37460f00",
        1289 => x"13060624",
        1290 => x"93060000",
        1291 => x"13050900",
        1292 => x"93050400",
        1293 => x"eff05fb5",
        1294 => x"37460f00",
        1295 => x"23a4a400",
        1296 => x"93050400",
        1297 => x"13050900",
        1298 => x"13060624",
        1299 => x"93060000",
        1300 => x"eff08ff0",
        1301 => x"8320c100",
        1302 => x"03248100",
        1303 => x"23a0a400",
        1304 => x"23a2b400",
        1305 => x"03290100",
        1306 => x"83244100",
        1307 => x"13050000",
        1308 => x"13010101",
        1309 => x"67800000",
        1310 => x"03a74188",
        1311 => x"b7870020",
        1312 => x"93870700",
        1313 => x"93060040",
        1314 => x"b387d740",
        1315 => x"630c0700",
        1316 => x"3305a700",
        1317 => x"63e2a702",
        1318 => x"23a2a188",
        1319 => x"13050700",
        1320 => x"67800000",
        1321 => x"93868189",
        1322 => x"13878189",
        1323 => x"23a2d188",
        1324 => x"3305a700",
        1325 => x"e3f2a7fe",
        1326 => x"130101ff",
        1327 => x"23261100",
        1328 => x"ef000032",
        1329 => x"8320c100",
        1330 => x"9307c000",
        1331 => x"2320f500",
        1332 => x"1307f0ff",
        1333 => x"13050700",
        1334 => x"13010101",
        1335 => x"67800000",
        1336 => x"130101f9",
        1337 => x"23248106",
        1338 => x"23229106",
        1339 => x"23261106",
        1340 => x"23202107",
        1341 => x"232e3105",
        1342 => x"232c4105",
        1343 => x"232a5105",
        1344 => x"23286105",
        1345 => x"23267105",
        1346 => x"23248105",
        1347 => x"23229105",
        1348 => x"2320a105",
        1349 => x"93040500",
        1350 => x"13840500",
        1351 => x"232c0100",
        1352 => x"232e0100",
        1353 => x"23200102",
        1354 => x"23220102",
        1355 => x"23240102",
        1356 => x"23260102",
        1357 => x"23280102",
        1358 => x"232a0102",
        1359 => x"232c0102",
        1360 => x"232e0102",
        1361 => x"97f2ffff",
        1362 => x"938282d3",
        1363 => x"73905230",
        1364 => x"93050004",
        1365 => x"1305101b",
        1366 => x"eff08f91",
        1367 => x"37877d01",
        1368 => x"b70700f0",
        1369 => x"1307f783",
        1370 => x"23a6e708",
        1371 => x"93061001",
        1372 => x"37170000",
        1373 => x"23a0d708",
        1374 => x"13077738",
        1375 => x"23a8e70a",
        1376 => x"37270000",
        1377 => x"1307f770",
        1378 => x"23a6e70a",
        1379 => x"23a0d70a",
        1380 => x"13078070",
        1381 => x"23a0e706",
        1382 => x"3707f900",
        1383 => x"13078700",
        1384 => x"23a0e704",
        1385 => x"93020008",
        1386 => x"73904230",
        1387 => x"b7220000",
        1388 => x"93828280",
        1389 => x"73900230",
        1390 => x"b7390000",
        1391 => x"138509e6",
        1392 => x"eff00f8e",
        1393 => x"63549002",
        1394 => x"1389f4ff",
        1395 => x"9304f0ff",
        1396 => x"03250400",
        1397 => x"1309f9ff",
        1398 => x"13044400",
        1399 => x"eff04f8c",
        1400 => x"138509e6",
        1401 => x"eff0cf8b",
        1402 => x"e31499fe",
        1403 => x"37350000",
        1404 => x"b7faeeee",
        1405 => x"130545e3",
        1406 => x"b7090010",
        1407 => x"37140000",
        1408 => x"1389faee",
        1409 => x"eff0cf89",
        1410 => x"373b0000",
        1411 => x"9389f9ff",
        1412 => x"938aeaee",
        1413 => x"130404e1",
        1414 => x"93040000",
        1415 => x"b71b0000",
        1416 => x"938b0b2c",
        1417 => x"130af000",
        1418 => x"93050000",
        1419 => x"13058100",
        1420 => x"ef008036",
        1421 => x"938bfbff",
        1422 => x"630a0502",
        1423 => x"e3960bfe",
        1424 => x"73001000",
        1425 => x"b70700f0",
        1426 => x"9306f00f",
        1427 => x"23a4d706",
        1428 => x"03a70704",
        1429 => x"93860704",
        1430 => x"13670730",
        1431 => x"23a0e704",
        1432 => x"93070009",
        1433 => x"23a4f600",
        1434 => x"6ff05ffb",
        1435 => x"032c8100",
        1436 => x"8325c100",
        1437 => x"13060400",
        1438 => x"9357cc01",
        1439 => x"13974500",
        1440 => x"b367f700",
        1441 => x"b3f73701",
        1442 => x"33773c01",
        1443 => x"13d5f541",
        1444 => x"13d88501",
        1445 => x"3307f700",
        1446 => x"33070701",
        1447 => x"9377d500",
        1448 => x"3307f700",
        1449 => x"33774703",
        1450 => x"937725ff",
        1451 => x"93860400",
        1452 => x"13050c00",
        1453 => x"3307f700",
        1454 => x"b307ec40",
        1455 => x"1357f741",
        1456 => x"3338fc00",
        1457 => x"3387e540",
        1458 => x"33070741",
        1459 => x"b3885703",
        1460 => x"33072703",
        1461 => x"33b82703",
        1462 => x"33071701",
        1463 => x"b3872703",
        1464 => x"33070701",
        1465 => x"1358f741",
        1466 => x"13783800",
        1467 => x"b307f800",
        1468 => x"33b80701",
        1469 => x"3307e800",
        1470 => x"1318e701",
        1471 => x"93d72700",
        1472 => x"b367f800",
        1473 => x"13582740",
        1474 => x"93184800",
        1475 => x"13d3c701",
        1476 => x"33e36800",
        1477 => x"33733301",
        1478 => x"b3f83701",
        1479 => x"135e8801",
        1480 => x"1357f741",
        1481 => x"b3886800",
        1482 => x"b388c801",
        1483 => x"1373d700",
        1484 => x"b3886800",
        1485 => x"b3f84803",
        1486 => x"137727ff",
        1487 => x"939c4700",
        1488 => x"b38cfc40",
        1489 => x"939c2c00",
        1490 => x"b30c9c41",
        1491 => x"b388e800",
        1492 => x"33871741",
        1493 => x"93d8f841",
        1494 => x"33b3e700",
        1495 => x"33081841",
        1496 => x"33086840",
        1497 => x"33082803",
        1498 => x"33035703",
        1499 => x"b3382703",
        1500 => x"33086800",
        1501 => x"33072703",
        1502 => x"33081801",
        1503 => x"9358f841",
        1504 => x"93f83800",
        1505 => x"3387e800",
        1506 => x"b3381701",
        1507 => x"b3880801",
        1508 => x"9398e801",
        1509 => x"13572700",
        1510 => x"33e7e800",
        1511 => x"13184700",
        1512 => x"3307e840",
        1513 => x"13172700",
        1514 => x"338de740",
        1515 => x"efe05ff3",
        1516 => x"83260101",
        1517 => x"13070500",
        1518 => x"13880c00",
        1519 => x"93070d00",
        1520 => x"13060c00",
        1521 => x"93054be6",
        1522 => x"13058101",
        1523 => x"ef00c015",
        1524 => x"13058101",
        1525 => x"efe0dfec",
        1526 => x"e3980be4",
        1527 => x"6ff05fe6",
        1528 => x"03a5c187",
        1529 => x"67800000",
        1530 => x"130101ff",
        1531 => x"23248100",
        1532 => x"23261100",
        1533 => x"93070000",
        1534 => x"13040500",
        1535 => x"63880700",
        1536 => x"93050000",
        1537 => x"97000000",
        1538 => x"e7000000",
        1539 => x"b7370000",
        1540 => x"03a547fc",
        1541 => x"83278502",
        1542 => x"63840700",
        1543 => x"e7800700",
        1544 => x"13050400",
        1545 => x"eff05fbc",
        1546 => x"130101ff",
        1547 => x"23248100",
        1548 => x"23229100",
        1549 => x"37340000",
        1550 => x"b7340000",
        1551 => x"938784fc",
        1552 => x"130484fc",
        1553 => x"3304f440",
        1554 => x"23202101",
        1555 => x"23261100",
        1556 => x"13542440",
        1557 => x"938484fc",
        1558 => x"13090000",
        1559 => x"63108904",
        1560 => x"b7340000",
        1561 => x"37340000",
        1562 => x"938784fc",
        1563 => x"130484fc",
        1564 => x"3304f440",
        1565 => x"13542440",
        1566 => x"938484fc",
        1567 => x"13090000",
        1568 => x"63188902",
        1569 => x"8320c100",
        1570 => x"03248100",
        1571 => x"83244100",
        1572 => x"03290100",
        1573 => x"13010101",
        1574 => x"67800000",
        1575 => x"83a70400",
        1576 => x"13091900",
        1577 => x"93844400",
        1578 => x"e7800700",
        1579 => x"6ff01ffb",
        1580 => x"83a70400",
        1581 => x"13091900",
        1582 => x"93844400",
        1583 => x"e7800700",
        1584 => x"6ff01ffc",
        1585 => x"130101f6",
        1586 => x"232af108",
        1587 => x"b7070080",
        1588 => x"93c7f7ff",
        1589 => x"232ef100",
        1590 => x"2328f100",
        1591 => x"b707ffff",
        1592 => x"2326d108",
        1593 => x"2324b100",
        1594 => x"232cb100",
        1595 => x"93878720",
        1596 => x"9306c108",
        1597 => x"93058100",
        1598 => x"232e1106",
        1599 => x"232af100",
        1600 => x"2328e108",
        1601 => x"232c0109",
        1602 => x"232e1109",
        1603 => x"2322d100",
        1604 => x"ef00c040",
        1605 => x"83278100",
        1606 => x"23800700",
        1607 => x"8320c107",
        1608 => x"1301010a",
        1609 => x"67800000",
        1610 => x"130101f6",
        1611 => x"232af108",
        1612 => x"b7070080",
        1613 => x"93c7f7ff",
        1614 => x"232ef100",
        1615 => x"2328f100",
        1616 => x"b707ffff",
        1617 => x"93878720",
        1618 => x"232af100",
        1619 => x"2324a100",
        1620 => x"232ca100",
        1621 => x"03a5c187",
        1622 => x"2324c108",
        1623 => x"2326d108",
        1624 => x"13860500",
        1625 => x"93068108",
        1626 => x"93058100",
        1627 => x"232e1106",
        1628 => x"2328e108",
        1629 => x"232c0109",
        1630 => x"232e1109",
        1631 => x"2322d100",
        1632 => x"ef00c039",
        1633 => x"83278100",
        1634 => x"23800700",
        1635 => x"8320c107",
        1636 => x"1301010a",
        1637 => x"67800000",
        1638 => x"13860500",
        1639 => x"93050500",
        1640 => x"03a5c187",
        1641 => x"6f004000",
        1642 => x"130101ff",
        1643 => x"23248100",
        1644 => x"23229100",
        1645 => x"13040500",
        1646 => x"13850500",
        1647 => x"93050600",
        1648 => x"23261100",
        1649 => x"23a40188",
        1650 => x"eff05fa2",
        1651 => x"9307f0ff",
        1652 => x"6318f500",
        1653 => x"83a78188",
        1654 => x"63840700",
        1655 => x"2320f400",
        1656 => x"8320c100",
        1657 => x"03248100",
        1658 => x"83244100",
        1659 => x"13010101",
        1660 => x"67800000",
        1661 => x"130101fe",
        1662 => x"23282101",
        1663 => x"03a98500",
        1664 => x"232c8100",
        1665 => x"23263101",
        1666 => x"23225101",
        1667 => x"23206101",
        1668 => x"232e1100",
        1669 => x"232a9100",
        1670 => x"23244101",
        1671 => x"83aa0500",
        1672 => x"13840500",
        1673 => x"130b0600",
        1674 => x"93890600",
        1675 => x"63ec2609",
        1676 => x"8397c500",
        1677 => x"13f70748",
        1678 => x"63040708",
        1679 => x"03274401",
        1680 => x"93043000",
        1681 => x"83a50501",
        1682 => x"b384e402",
        1683 => x"13072000",
        1684 => x"b38aba40",
        1685 => x"130a0500",
        1686 => x"b3c4e402",
        1687 => x"13871600",
        1688 => x"33075701",
        1689 => x"63f4e400",
        1690 => x"93040700",
        1691 => x"93f70740",
        1692 => x"6386070a",
        1693 => x"93850400",
        1694 => x"13050a00",
        1695 => x"ef001067",
        1696 => x"13090500",
        1697 => x"630c050a",
        1698 => x"83250401",
        1699 => x"13860a00",
        1700 => x"eff0df8d",
        1701 => x"8357c400",
        1702 => x"93f7f7b7",
        1703 => x"93e70708",
        1704 => x"2316f400",
        1705 => x"23282401",
        1706 => x"232a9400",
        1707 => x"33095901",
        1708 => x"b3845441",
        1709 => x"23202401",
        1710 => x"23249400",
        1711 => x"13890900",
        1712 => x"63f42901",
        1713 => x"13890900",
        1714 => x"03250400",
        1715 => x"13060900",
        1716 => x"93050b00",
        1717 => x"eff09f8d",
        1718 => x"83278400",
        1719 => x"13050000",
        1720 => x"b3872741",
        1721 => x"2324f400",
        1722 => x"83270400",
        1723 => x"b3872701",
        1724 => x"2320f400",
        1725 => x"8320c101",
        1726 => x"03248101",
        1727 => x"83244101",
        1728 => x"03290101",
        1729 => x"8329c100",
        1730 => x"032a8100",
        1731 => x"832a4100",
        1732 => x"032b0100",
        1733 => x"13010102",
        1734 => x"67800000",
        1735 => x"13860400",
        1736 => x"13050a00",
        1737 => x"ef001071",
        1738 => x"13090500",
        1739 => x"e31c05f6",
        1740 => x"83250401",
        1741 => x"13050a00",
        1742 => x"ef00d04b",
        1743 => x"9307c000",
        1744 => x"2320fa00",
        1745 => x"8357c400",
        1746 => x"1305f0ff",
        1747 => x"93e70704",
        1748 => x"2316f400",
        1749 => x"6ff01ffa",
        1750 => x"83278600",
        1751 => x"130101fd",
        1752 => x"232e3101",
        1753 => x"23286101",
        1754 => x"23261102",
        1755 => x"23248102",
        1756 => x"23229102",
        1757 => x"23202103",
        1758 => x"232c4101",
        1759 => x"232a5101",
        1760 => x"23267101",
        1761 => x"23248101",
        1762 => x"23229101",
        1763 => x"2320a101",
        1764 => x"032b0600",
        1765 => x"93090600",
        1766 => x"63940712",
        1767 => x"13050000",
        1768 => x"8320c102",
        1769 => x"03248102",
        1770 => x"23a20900",
        1771 => x"83244102",
        1772 => x"03290102",
        1773 => x"8329c101",
        1774 => x"032a8101",
        1775 => x"832a4101",
        1776 => x"032b0101",
        1777 => x"832bc100",
        1778 => x"032c8100",
        1779 => x"832c4100",
        1780 => x"032d0100",
        1781 => x"13010103",
        1782 => x"67800000",
        1783 => x"832b0b00",
        1784 => x"032d4b00",
        1785 => x"130b8b00",
        1786 => x"03298400",
        1787 => x"832a0400",
        1788 => x"e3060dfe",
        1789 => x"63642d09",
        1790 => x"8317c400",
        1791 => x"13f70748",
        1792 => x"630e0706",
        1793 => x"83244401",
        1794 => x"83250401",
        1795 => x"b3049c02",
        1796 => x"b38aba40",
        1797 => x"13871a00",
        1798 => x"3307a701",
        1799 => x"b3c49403",
        1800 => x"63f4e400",
        1801 => x"93040700",
        1802 => x"93f70740",
        1803 => x"6388070a",
        1804 => x"93850400",
        1805 => x"13050a00",
        1806 => x"ef00504b",
        1807 => x"13090500",
        1808 => x"630e050a",
        1809 => x"83250401",
        1810 => x"13860a00",
        1811 => x"eff00ff2",
        1812 => x"8357c400",
        1813 => x"93f7f7b7",
        1814 => x"93e70708",
        1815 => x"2316f400",
        1816 => x"23282401",
        1817 => x"232a9400",
        1818 => x"33095901",
        1819 => x"b3845441",
        1820 => x"23202401",
        1821 => x"23249400",
        1822 => x"13090d00",
        1823 => x"63742d01",
        1824 => x"13090d00",
        1825 => x"03250400",
        1826 => x"13060900",
        1827 => x"93850b00",
        1828 => x"eff0cff1",
        1829 => x"83278400",
        1830 => x"b3872741",
        1831 => x"2324f400",
        1832 => x"83270400",
        1833 => x"b3872701",
        1834 => x"2320f400",
        1835 => x"83a78900",
        1836 => x"b387a741",
        1837 => x"23a4f900",
        1838 => x"e39207f2",
        1839 => x"6ff01fee",
        1840 => x"130a0500",
        1841 => x"13840500",
        1842 => x"930b0000",
        1843 => x"130d0000",
        1844 => x"130c3000",
        1845 => x"930c2000",
        1846 => x"6ff01ff1",
        1847 => x"13860400",
        1848 => x"13050a00",
        1849 => x"ef001055",
        1850 => x"13090500",
        1851 => x"e31a05f6",
        1852 => x"83250401",
        1853 => x"13050a00",
        1854 => x"ef00d02f",
        1855 => x"9307c000",
        1856 => x"2320fa00",
        1857 => x"8357c400",
        1858 => x"1305f0ff",
        1859 => x"93e70704",
        1860 => x"2316f400",
        1861 => x"23a40900",
        1862 => x"6ff09fe8",
        1863 => x"83d7c500",
        1864 => x"130101f5",
        1865 => x"2324810a",
        1866 => x"2322910a",
        1867 => x"2320210b",
        1868 => x"232c4109",
        1869 => x"2326110a",
        1870 => x"232e3109",
        1871 => x"232a5109",
        1872 => x"23286109",
        1873 => x"23267109",
        1874 => x"23248109",
        1875 => x"23229109",
        1876 => x"2320a109",
        1877 => x"232eb107",
        1878 => x"93f70708",
        1879 => x"130a0500",
        1880 => x"13890500",
        1881 => x"93040600",
        1882 => x"13840600",
        1883 => x"63880706",
        1884 => x"83a70501",
        1885 => x"63940706",
        1886 => x"93050004",
        1887 => x"ef001037",
        1888 => x"2320a900",
        1889 => x"2328a900",
        1890 => x"63160504",
        1891 => x"9307c000",
        1892 => x"2320fa00",
        1893 => x"1305f0ff",
        1894 => x"8320c10a",
        1895 => x"0324810a",
        1896 => x"8324410a",
        1897 => x"0329010a",
        1898 => x"8329c109",
        1899 => x"032a8109",
        1900 => x"832a4109",
        1901 => x"032b0109",
        1902 => x"832bc108",
        1903 => x"032c8108",
        1904 => x"832c4108",
        1905 => x"032d0108",
        1906 => x"832dc107",
        1907 => x"1301010b",
        1908 => x"67800000",
        1909 => x"93070004",
        1910 => x"232af900",
        1911 => x"93070002",
        1912 => x"a304f102",
        1913 => x"93070003",
        1914 => x"23220102",
        1915 => x"2305f102",
        1916 => x"23268100",
        1917 => x"930c5002",
        1918 => x"373b0000",
        1919 => x"b73b0000",
        1920 => x"373d0000",
        1921 => x"372c0000",
        1922 => x"930a0000",
        1923 => x"13840400",
        1924 => x"83470400",
        1925 => x"63840700",
        1926 => x"639c970d",
        1927 => x"b30d9440",
        1928 => x"63069402",
        1929 => x"93860d00",
        1930 => x"13860400",
        1931 => x"93050900",
        1932 => x"13050a00",
        1933 => x"eff01fbc",
        1934 => x"9307f0ff",
        1935 => x"6304f524",
        1936 => x"83274102",
        1937 => x"b387b701",
        1938 => x"2322f102",
        1939 => x"83470400",
        1940 => x"638a0722",
        1941 => x"9307f0ff",
        1942 => x"93041400",
        1943 => x"23280100",
        1944 => x"232e0100",
        1945 => x"232af100",
        1946 => x"232c0100",
        1947 => x"a3090104",
        1948 => x"23240106",
        1949 => x"930d1000",
        1950 => x"83c50400",
        1951 => x"13065000",
        1952 => x"13050bf3",
        1953 => x"ef00d014",
        1954 => x"83270101",
        1955 => x"13841400",
        1956 => x"63140506",
        1957 => x"13f70701",
        1958 => x"63060700",
        1959 => x"13070002",
        1960 => x"a309e104",
        1961 => x"13f78700",
        1962 => x"63060700",
        1963 => x"1307b002",
        1964 => x"a309e104",
        1965 => x"83c60400",
        1966 => x"1307a002",
        1967 => x"638ce604",
        1968 => x"8327c101",
        1969 => x"13840400",
        1970 => x"93060000",
        1971 => x"13069000",
        1972 => x"1305a000",
        1973 => x"03470400",
        1974 => x"93051400",
        1975 => x"130707fd",
        1976 => x"637ee608",
        1977 => x"63840604",
        1978 => x"232ef100",
        1979 => x"6f000004",
        1980 => x"13041400",
        1981 => x"6ff0dff1",
        1982 => x"13070bf3",
        1983 => x"3305e540",
        1984 => x"3395ad00",
        1985 => x"b3e7a700",
        1986 => x"2328f100",
        1987 => x"93040400",
        1988 => x"6ff09ff6",
        1989 => x"0327c100",
        1990 => x"93064700",
        1991 => x"03270700",
        1992 => x"2326d100",
        1993 => x"63420704",
        1994 => x"232ee100",
        1995 => x"03470400",
        1996 => x"9307e002",
        1997 => x"6314f708",
        1998 => x"03471400",
        1999 => x"9307a002",
        2000 => x"6318f704",
        2001 => x"8327c100",
        2002 => x"13042400",
        2003 => x"13874700",
        2004 => x"83a70700",
        2005 => x"2326e100",
        2006 => x"63d40700",
        2007 => x"9307f0ff",
        2008 => x"232af100",
        2009 => x"6f008005",
        2010 => x"3307e040",
        2011 => x"93e72700",
        2012 => x"232ee100",
        2013 => x"2328f100",
        2014 => x"6ff05ffb",
        2015 => x"b387a702",
        2016 => x"13840500",
        2017 => x"93061000",
        2018 => x"b387e700",
        2019 => x"6ff09ff4",
        2020 => x"13041400",
        2021 => x"232a0100",
        2022 => x"93060000",
        2023 => x"93070000",
        2024 => x"13069000",
        2025 => x"1305a000",
        2026 => x"03470400",
        2027 => x"93051400",
        2028 => x"130707fd",
        2029 => x"6372e608",
        2030 => x"e39406fa",
        2031 => x"83450400",
        2032 => x"13063000",
        2033 => x"13858bf3",
        2034 => x"ef009000",
        2035 => x"63020502",
        2036 => x"93878bf3",
        2037 => x"3305f540",
        2038 => x"83270101",
        2039 => x"13070004",
        2040 => x"3317a700",
        2041 => x"b3e7e700",
        2042 => x"13041400",
        2043 => x"2328f100",
        2044 => x"83450400",
        2045 => x"13066000",
        2046 => x"1305cdf3",
        2047 => x"93041400",
        2048 => x"2304b102",
        2049 => x"ef00c07c",
        2050 => x"63080508",
        2051 => x"63980a04",
        2052 => x"03270101",
        2053 => x"8327c100",
        2054 => x"13770710",
        2055 => x"63080702",
        2056 => x"93874700",
        2057 => x"2326f100",
        2058 => x"83274102",
        2059 => x"b3873701",
        2060 => x"2322f102",
        2061 => x"6ff09fdd",
        2062 => x"b387a702",
        2063 => x"13840500",
        2064 => x"93061000",
        2065 => x"b387e700",
        2066 => x"6ff01ff6",
        2067 => x"93877700",
        2068 => x"93f787ff",
        2069 => x"93878700",
        2070 => x"6ff0dffc",
        2071 => x"1307c100",
        2072 => x"93064c9f",
        2073 => x"13060900",
        2074 => x"93050101",
        2075 => x"13050a00",
        2076 => x"97000000",
        2077 => x"e7000000",
        2078 => x"9307f0ff",
        2079 => x"93090500",
        2080 => x"e314f5fa",
        2081 => x"8357c900",
        2082 => x"93f70704",
        2083 => x"e39407d0",
        2084 => x"03254102",
        2085 => x"6ff05fd0",
        2086 => x"1307c100",
        2087 => x"93064c9f",
        2088 => x"13060900",
        2089 => x"93050101",
        2090 => x"13050a00",
        2091 => x"ef00801b",
        2092 => x"6ff09ffc",
        2093 => x"130101fd",
        2094 => x"232a5101",
        2095 => x"83a70501",
        2096 => x"930a0700",
        2097 => x"03a78500",
        2098 => x"23248102",
        2099 => x"23202103",
        2100 => x"232e3101",
        2101 => x"232c4101",
        2102 => x"23261102",
        2103 => x"23229102",
        2104 => x"23286101",
        2105 => x"23267101",
        2106 => x"93090500",
        2107 => x"13840500",
        2108 => x"13090600",
        2109 => x"138a0600",
        2110 => x"63d4e700",
        2111 => x"93070700",
        2112 => x"2320f900",
        2113 => x"03473404",
        2114 => x"63060700",
        2115 => x"93871700",
        2116 => x"2320f900",
        2117 => x"83270400",
        2118 => x"93f70702",
        2119 => x"63880700",
        2120 => x"83270900",
        2121 => x"93872700",
        2122 => x"2320f900",
        2123 => x"83240400",
        2124 => x"93f46400",
        2125 => x"639e0400",
        2126 => x"130b9401",
        2127 => x"930bf0ff",
        2128 => x"8327c400",
        2129 => x"03270900",
        2130 => x"b387e740",
        2131 => x"63c2f408",
        2132 => x"83473404",
        2133 => x"b336f000",
        2134 => x"83270400",
        2135 => x"93f70702",
        2136 => x"6390070c",
        2137 => x"13063404",
        2138 => x"93050a00",
        2139 => x"13850900",
        2140 => x"e7800a00",
        2141 => x"9307f0ff",
        2142 => x"6308f506",
        2143 => x"83270400",
        2144 => x"13074000",
        2145 => x"93040000",
        2146 => x"93f76700",
        2147 => x"639ce700",
        2148 => x"8324c400",
        2149 => x"83270900",
        2150 => x"b384f440",
        2151 => x"63d40400",
        2152 => x"93040000",
        2153 => x"83278400",
        2154 => x"03270401",
        2155 => x"6356f700",
        2156 => x"b387e740",
        2157 => x"b384f400",
        2158 => x"13090000",
        2159 => x"1304a401",
        2160 => x"130bf0ff",
        2161 => x"63902409",
        2162 => x"13050000",
        2163 => x"6f000002",
        2164 => x"93061000",
        2165 => x"13060b00",
        2166 => x"93050a00",
        2167 => x"13850900",
        2168 => x"e7800a00",
        2169 => x"631a7503",
        2170 => x"1305f0ff",
        2171 => x"8320c102",
        2172 => x"03248102",
        2173 => x"83244102",
        2174 => x"03290102",
        2175 => x"8329c101",
        2176 => x"032a8101",
        2177 => x"832a4101",
        2178 => x"032b0101",
        2179 => x"832bc100",
        2180 => x"13010103",
        2181 => x"67800000",
        2182 => x"93841400",
        2183 => x"6ff05ff2",
        2184 => x"3307d400",
        2185 => x"13060003",
        2186 => x"a301c704",
        2187 => x"03475404",
        2188 => x"93871600",
        2189 => x"b307f400",
        2190 => x"93862600",
        2191 => x"a381e704",
        2192 => x"6ff05ff2",
        2193 => x"93061000",
        2194 => x"13060400",
        2195 => x"93050a00",
        2196 => x"13850900",
        2197 => x"e7800a00",
        2198 => x"e30865f9",
        2199 => x"13091900",
        2200 => x"6ff05ff6",
        2201 => x"130101fd",
        2202 => x"23248102",
        2203 => x"23229102",
        2204 => x"23202103",
        2205 => x"232e3101",
        2206 => x"23261102",
        2207 => x"232c4101",
        2208 => x"232a5101",
        2209 => x"23286101",
        2210 => x"83c88501",
        2211 => x"93078007",
        2212 => x"93040500",
        2213 => x"13840500",
        2214 => x"13090600",
        2215 => x"93890600",
        2216 => x"63ee1701",
        2217 => x"93072006",
        2218 => x"93863504",
        2219 => x"63ee1701",
        2220 => x"638a082a",
        2221 => x"93078005",
        2222 => x"638af820",
        2223 => x"930a2404",
        2224 => x"23011405",
        2225 => x"6f004004",
        2226 => x"9387d8f9",
        2227 => x"93f7f70f",
        2228 => x"13065001",
        2229 => x"e364f6fe",
        2230 => x"37360000",
        2231 => x"93972700",
        2232 => x"1306c6f6",
        2233 => x"b387c700",
        2234 => x"83a70700",
        2235 => x"67800700",
        2236 => x"83270700",
        2237 => x"938a2504",
        2238 => x"93864700",
        2239 => x"83a70700",
        2240 => x"2320d700",
        2241 => x"2381f504",
        2242 => x"93071000",
        2243 => x"6f004029",
        2244 => x"03a60500",
        2245 => x"83270700",
        2246 => x"13750608",
        2247 => x"93854700",
        2248 => x"630e0504",
        2249 => x"83a70700",
        2250 => x"2320b700",
        2251 => x"37370000",
        2252 => x"83254400",
        2253 => x"130847f4",
        2254 => x"63d2071e",
        2255 => x"1307d002",
        2256 => x"a301e404",
        2257 => x"2324b400",
        2258 => x"63d80504",
        2259 => x"b307f040",
        2260 => x"1307a000",
        2261 => x"938a0600",
        2262 => x"33f6e702",
        2263 => x"938afaff",
        2264 => x"3306c800",
        2265 => x"03460600",
        2266 => x"2380ca00",
        2267 => x"13860700",
        2268 => x"b3d7e702",
        2269 => x"e372e6fe",
        2270 => x"6f008009",
        2271 => x"83a70700",
        2272 => x"13750604",
        2273 => x"2320b700",
        2274 => x"e30205fa",
        2275 => x"93970701",
        2276 => x"93d70741",
        2277 => x"6ff09ff9",
        2278 => x"1376b6ff",
        2279 => x"2320c400",
        2280 => x"6ff0dffa",
        2281 => x"03a60500",
        2282 => x"83270700",
        2283 => x"13750608",
        2284 => x"93854700",
        2285 => x"63080500",
        2286 => x"2320b700",
        2287 => x"83a70700",
        2288 => x"6f004001",
        2289 => x"13760604",
        2290 => x"2320b700",
        2291 => x"e30806fe",
        2292 => x"83d70700",
        2293 => x"37380000",
        2294 => x"1307f006",
        2295 => x"130848f4",
        2296 => x"639ae812",
        2297 => x"13078000",
        2298 => x"a3010404",
        2299 => x"03264400",
        2300 => x"2324c400",
        2301 => x"e34006f6",
        2302 => x"83250400",
        2303 => x"93f5b5ff",
        2304 => x"2320b400",
        2305 => x"e39807f4",
        2306 => x"938a0600",
        2307 => x"e31406f4",
        2308 => x"93078000",
        2309 => x"6314f702",
        2310 => x"83270400",
        2311 => x"93f71700",
        2312 => x"638e0700",
        2313 => x"03274400",
        2314 => x"83270401",
        2315 => x"63c8e700",
        2316 => x"93070003",
        2317 => x"a38ffafe",
        2318 => x"938afaff",
        2319 => x"b3865641",
        2320 => x"2328d400",
        2321 => x"13870900",
        2322 => x"93060900",
        2323 => x"1306c100",
        2324 => x"93050400",
        2325 => x"13850400",
        2326 => x"eff0dfc5",
        2327 => x"130af0ff",
        2328 => x"63164515",
        2329 => x"1305f0ff",
        2330 => x"8320c102",
        2331 => x"03248102",
        2332 => x"83244102",
        2333 => x"03290102",
        2334 => x"8329c101",
        2335 => x"032a8101",
        2336 => x"832a4101",
        2337 => x"032b0101",
        2338 => x"13010103",
        2339 => x"67800000",
        2340 => x"83a70500",
        2341 => x"93e70702",
        2342 => x"23a0f500",
        2343 => x"37380000",
        2344 => x"93088007",
        2345 => x"130888f5",
        2346 => x"03260400",
        2347 => x"a3021405",
        2348 => x"83270700",
        2349 => x"13750608",
        2350 => x"93854700",
        2351 => x"630e0500",
        2352 => x"2320b700",
        2353 => x"83a70700",
        2354 => x"6f000002",
        2355 => x"37380000",
        2356 => x"130848f4",
        2357 => x"6ff05ffd",
        2358 => x"13750604",
        2359 => x"2320b700",
        2360 => x"e30205fe",
        2361 => x"83d70700",
        2362 => x"13771600",
        2363 => x"63060700",
        2364 => x"13660602",
        2365 => x"2320c400",
        2366 => x"63860700",
        2367 => x"13070001",
        2368 => x"6ff09fee",
        2369 => x"03270400",
        2370 => x"1377f7fd",
        2371 => x"2320e400",
        2372 => x"6ff0dffe",
        2373 => x"1307a000",
        2374 => x"6ff01fed",
        2375 => x"130847f4",
        2376 => x"1307a000",
        2377 => x"6ff09fec",
        2378 => x"03a60500",
        2379 => x"83270700",
        2380 => x"83a54501",
        2381 => x"13780608",
        2382 => x"13854700",
        2383 => x"630a0800",
        2384 => x"2320a700",
        2385 => x"83a70700",
        2386 => x"23a0b700",
        2387 => x"6f008001",
        2388 => x"2320a700",
        2389 => x"13760604",
        2390 => x"83a70700",
        2391 => x"e30606fe",
        2392 => x"2390b700",
        2393 => x"23280400",
        2394 => x"938a0600",
        2395 => x"6ff09fed",
        2396 => x"83270700",
        2397 => x"03a64500",
        2398 => x"93050000",
        2399 => x"93864700",
        2400 => x"2320d700",
        2401 => x"83aa0700",
        2402 => x"13850a00",
        2403 => x"ef004024",
        2404 => x"63060500",
        2405 => x"33055541",
        2406 => x"2322a400",
        2407 => x"83274400",
        2408 => x"2328f400",
        2409 => x"a3010404",
        2410 => x"6ff0dfe9",
        2411 => x"83260401",
        2412 => x"13860a00",
        2413 => x"93050900",
        2414 => x"13850400",
        2415 => x"e7800900",
        2416 => x"e30245eb",
        2417 => x"83270400",
        2418 => x"93f72700",
        2419 => x"63940704",
        2420 => x"8327c100",
        2421 => x"0325c400",
        2422 => x"e358f5e8",
        2423 => x"13850700",
        2424 => x"6ff09fe8",
        2425 => x"93061000",
        2426 => x"13860a00",
        2427 => x"93050900",
        2428 => x"13850400",
        2429 => x"e7800900",
        2430 => x"e30665e7",
        2431 => x"130a1a00",
        2432 => x"8327c400",
        2433 => x"0327c100",
        2434 => x"b387e740",
        2435 => x"e34cfafc",
        2436 => x"6ff01ffc",
        2437 => x"130a0000",
        2438 => x"930a9401",
        2439 => x"130bf0ff",
        2440 => x"6ff01ffe",
        2441 => x"130101ff",
        2442 => x"23248100",
        2443 => x"13840500",
        2444 => x"83a50500",
        2445 => x"23229100",
        2446 => x"23261100",
        2447 => x"93040500",
        2448 => x"63840500",
        2449 => x"eff01ffe",
        2450 => x"93050400",
        2451 => x"03248100",
        2452 => x"8320c100",
        2453 => x"13850400",
        2454 => x"83244100",
        2455 => x"13010101",
        2456 => x"6f004019",
        2457 => x"83a7c187",
        2458 => x"6382a716",
        2459 => x"83274502",
        2460 => x"130101fe",
        2461 => x"232c8100",
        2462 => x"232e1100",
        2463 => x"232a9100",
        2464 => x"23282101",
        2465 => x"23263101",
        2466 => x"13040500",
        2467 => x"638a0704",
        2468 => x"83a7c700",
        2469 => x"638c0702",
        2470 => x"93040000",
        2471 => x"13090008",
        2472 => x"83274402",
        2473 => x"83a7c700",
        2474 => x"b3879700",
        2475 => x"83a50700",
        2476 => x"6396050e",
        2477 => x"93844400",
        2478 => x"e39424ff",
        2479 => x"83274402",
        2480 => x"13050400",
        2481 => x"83a5c700",
        2482 => x"ef00c012",
        2483 => x"83274402",
        2484 => x"83a50700",
        2485 => x"63860500",
        2486 => x"13050400",
        2487 => x"ef008011",
        2488 => x"83254401",
        2489 => x"63860500",
        2490 => x"13050400",
        2491 => x"ef008010",
        2492 => x"83254402",
        2493 => x"63860500",
        2494 => x"13050400",
        2495 => x"ef00800f",
        2496 => x"83258403",
        2497 => x"63860500",
        2498 => x"13050400",
        2499 => x"ef00800e",
        2500 => x"8325c403",
        2501 => x"63860500",
        2502 => x"13050400",
        2503 => x"ef00800d",
        2504 => x"83250404",
        2505 => x"63860500",
        2506 => x"13050400",
        2507 => x"ef00800c",
        2508 => x"8325c405",
        2509 => x"63860500",
        2510 => x"13050400",
        2511 => x"ef00800b",
        2512 => x"83258405",
        2513 => x"63860500",
        2514 => x"13050400",
        2515 => x"ef00800a",
        2516 => x"83254403",
        2517 => x"63860500",
        2518 => x"13050400",
        2519 => x"ef008009",
        2520 => x"83278401",
        2521 => x"63860704",
        2522 => x"83278402",
        2523 => x"13050400",
        2524 => x"e7800700",
        2525 => x"83258404",
        2526 => x"638c0502",
        2527 => x"13050400",
        2528 => x"03248101",
        2529 => x"8320c101",
        2530 => x"83244101",
        2531 => x"03290101",
        2532 => x"8329c100",
        2533 => x"13010102",
        2534 => x"6ff0dfe8",
        2535 => x"83a90500",
        2536 => x"13050400",
        2537 => x"ef000005",
        2538 => x"93850900",
        2539 => x"6ff05ff0",
        2540 => x"8320c101",
        2541 => x"03248101",
        2542 => x"83244101",
        2543 => x"03290101",
        2544 => x"8329c100",
        2545 => x"13010102",
        2546 => x"67800000",
        2547 => x"67800000",
        2548 => x"93f5f50f",
        2549 => x"3306c500",
        2550 => x"6316c500",
        2551 => x"13050000",
        2552 => x"67800000",
        2553 => x"83470500",
        2554 => x"e38cb7fe",
        2555 => x"13051500",
        2556 => x"6ff09ffe",
        2557 => x"638a050e",
        2558 => x"83a7c5ff",
        2559 => x"130101fe",
        2560 => x"232c8100",
        2561 => x"232e1100",
        2562 => x"1384c5ff",
        2563 => x"63d40700",
        2564 => x"3304f400",
        2565 => x"2326a100",
        2566 => x"ef008033",
        2567 => x"83a70189",
        2568 => x"0325c100",
        2569 => x"639e0700",
        2570 => x"23220400",
        2571 => x"23a88188",
        2572 => x"03248101",
        2573 => x"8320c101",
        2574 => x"13010102",
        2575 => x"6f008031",
        2576 => x"6374f402",
        2577 => x"03260400",
        2578 => x"b306c400",
        2579 => x"639ad700",
        2580 => x"83a60700",
        2581 => x"83a74700",
        2582 => x"b386c600",
        2583 => x"2320d400",
        2584 => x"2322f400",
        2585 => x"6ff09ffc",
        2586 => x"13870700",
        2587 => x"83a74700",
        2588 => x"63840700",
        2589 => x"e37af4fe",
        2590 => x"83260700",
        2591 => x"3306d700",
        2592 => x"63188602",
        2593 => x"03260400",
        2594 => x"b386c600",
        2595 => x"2320d700",
        2596 => x"3306d700",
        2597 => x"e39ec7f8",
        2598 => x"03a60700",
        2599 => x"83a74700",
        2600 => x"b306d600",
        2601 => x"2320d700",
        2602 => x"2322f700",
        2603 => x"6ff05ff8",
        2604 => x"6378c400",
        2605 => x"9307c000",
        2606 => x"2320f500",
        2607 => x"6ff05ff7",
        2608 => x"03260400",
        2609 => x"b306c400",
        2610 => x"639ad700",
        2611 => x"83a60700",
        2612 => x"83a74700",
        2613 => x"b386c600",
        2614 => x"2320d400",
        2615 => x"2322f400",
        2616 => x"23228700",
        2617 => x"6ff0dff4",
        2618 => x"67800000",
        2619 => x"130101fe",
        2620 => x"232a9100",
        2621 => x"93843500",
        2622 => x"93f4c4ff",
        2623 => x"23282101",
        2624 => x"232e1100",
        2625 => x"232c8100",
        2626 => x"23263101",
        2627 => x"93848400",
        2628 => x"9307c000",
        2629 => x"13090500",
        2630 => x"63f0f406",
        2631 => x"9304c000",
        2632 => x"63eeb404",
        2633 => x"13050900",
        2634 => x"ef008022",
        2635 => x"03a70189",
        2636 => x"13040700",
        2637 => x"63180406",
        2638 => x"83a7c188",
        2639 => x"639a0700",
        2640 => x"93050000",
        2641 => x"13050900",
        2642 => x"ef00001c",
        2643 => x"23a6a188",
        2644 => x"93850400",
        2645 => x"13050900",
        2646 => x"ef00001b",
        2647 => x"9309f0ff",
        2648 => x"631a350b",
        2649 => x"9307c000",
        2650 => x"2320f900",
        2651 => x"13050900",
        2652 => x"ef00401e",
        2653 => x"6f000001",
        2654 => x"e3d404fa",
        2655 => x"9307c000",
        2656 => x"2320f900",
        2657 => x"13050000",
        2658 => x"8320c101",
        2659 => x"03248101",
        2660 => x"83244101",
        2661 => x"03290101",
        2662 => x"8329c100",
        2663 => x"13010102",
        2664 => x"67800000",
        2665 => x"83270400",
        2666 => x"b3879740",
        2667 => x"63ce0704",
        2668 => x"1306b000",
        2669 => x"637af600",
        2670 => x"2320f400",
        2671 => x"3304f400",
        2672 => x"23209400",
        2673 => x"6f000001",
        2674 => x"83274400",
        2675 => x"631a8702",
        2676 => x"23a8f188",
        2677 => x"13050900",
        2678 => x"ef00c017",
        2679 => x"1305b400",
        2680 => x"93074400",
        2681 => x"137585ff",
        2682 => x"3307f540",
        2683 => x"e30ef5f8",
        2684 => x"3304e400",
        2685 => x"b387a740",
        2686 => x"2320f400",
        2687 => x"6ff0dff8",
        2688 => x"2322f700",
        2689 => x"6ff01ffd",
        2690 => x"13070400",
        2691 => x"03244400",
        2692 => x"6ff05ff2",
        2693 => x"13043500",
        2694 => x"1374c4ff",
        2695 => x"e30285fa",
        2696 => x"b305a440",
        2697 => x"13050900",
        2698 => x"ef00000e",
        2699 => x"e31a35f9",
        2700 => x"6ff05ff3",
        2701 => x"130101fe",
        2702 => x"232c8100",
        2703 => x"232e1100",
        2704 => x"232a9100",
        2705 => x"23282101",
        2706 => x"23263101",
        2707 => x"23244101",
        2708 => x"13040600",
        2709 => x"63940502",
        2710 => x"03248101",
        2711 => x"8320c101",
        2712 => x"83244101",
        2713 => x"03290101",
        2714 => x"8329c100",
        2715 => x"032a8100",
        2716 => x"93050600",
        2717 => x"13010102",
        2718 => x"6ff05fe7",
        2719 => x"63180602",
        2720 => x"eff05fd7",
        2721 => x"93040000",
        2722 => x"8320c101",
        2723 => x"03248101",
        2724 => x"03290101",
        2725 => x"8329c100",
        2726 => x"032a8100",
        2727 => x"13850400",
        2728 => x"83244101",
        2729 => x"13010102",
        2730 => x"67800000",
        2731 => x"130a0500",
        2732 => x"93840500",
        2733 => x"ef00400a",
        2734 => x"13090500",
        2735 => x"63668500",
        2736 => x"93571500",
        2737 => x"e3e287fc",
        2738 => x"93050400",
        2739 => x"13050a00",
        2740 => x"eff0dfe1",
        2741 => x"93090500",
        2742 => x"e30605fa",
        2743 => x"13060400",
        2744 => x"63748900",
        2745 => x"13060900",
        2746 => x"93850400",
        2747 => x"13850900",
        2748 => x"efe0df87",
        2749 => x"93850400",
        2750 => x"13050a00",
        2751 => x"eff09fcf",
        2752 => x"93840900",
        2753 => x"6ff05ff8",
        2754 => x"130101ff",
        2755 => x"23248100",
        2756 => x"23229100",
        2757 => x"13040500",
        2758 => x"13850500",
        2759 => x"23261100",
        2760 => x"23a40188",
        2761 => x"efe05f95",
        2762 => x"9307f0ff",
        2763 => x"6318f500",
        2764 => x"83a78188",
        2765 => x"63840700",
        2766 => x"2320f400",
        2767 => x"8320c100",
        2768 => x"03248100",
        2769 => x"83244100",
        2770 => x"13010101",
        2771 => x"67800000",
        2772 => x"67800000",
        2773 => x"67800000",
        2774 => x"83a7c5ff",
        2775 => x"1385c7ff",
        2776 => x"63d80700",
        2777 => x"b385a500",
        2778 => x"83a70500",
        2779 => x"3305f500",
        2780 => x"67800000",
        2781 => x"10000000",
        2782 => x"00000000",
        2783 => x"037a5200",
        2784 => x"017c0101",
        2785 => x"1b0d0200",
        2786 => x"10000000",
        2787 => x"18000000",
        2788 => x"50dbffff",
        2789 => x"78040000",
        2790 => x"00000000",
        2791 => x"10000000",
        2792 => x"00000000",
        2793 => x"037a5200",
        2794 => x"017c0101",
        2795 => x"1b0d0200",
        2796 => x"10000000",
        2797 => x"18000000",
        2798 => x"a0dfffff",
        2799 => x"30040000",
        2800 => x"00000000",
        2801 => x"10000000",
        2802 => x"00000000",
        2803 => x"037a5200",
        2804 => x"017c0101",
        2805 => x"1b0d0200",
        2806 => x"10000000",
        2807 => x"18000000",
        2808 => x"a8e3ffff",
        2809 => x"e4030000",
        2810 => x"00000000",
        2811 => x"30313233",
        2812 => x"34353637",
        2813 => x"38396162",
        2814 => x"63646566",
        2815 => x"00000000",
        2816 => x"44040000",
        2817 => x"20040000",
        2818 => x"38040000",
        2819 => x"2c040000",
        2820 => x"74030000",
        2821 => x"74030000",
        2822 => x"74030000",
        2823 => x"88040000",
        2824 => x"74030000",
        2825 => x"74030000",
        2826 => x"74030000",
        2827 => x"74030000",
        2828 => x"74030000",
        2829 => x"74030000",
        2830 => x"74030000",
        2831 => x"50040000",
        2832 => x"ec040000",
        2833 => x"a4040000",
        2834 => x"a4040000",
        2835 => x"a4040000",
        2836 => x"a4040000",
        2837 => x"e0040000",
        2838 => x"2c050000",
        2839 => x"04050000",
        2840 => x"a4040000",
        2841 => x"a4040000",
        2842 => x"a4040000",
        2843 => x"a4040000",
        2844 => x"a4040000",
        2845 => x"a4040000",
        2846 => x"a4040000",
        2847 => x"a4040000",
        2848 => x"a4040000",
        2849 => x"a4040000",
        2850 => x"a4040000",
        2851 => x"a4040000",
        2852 => x"a4040000",
        2853 => x"a4040000",
        2854 => x"cc040000",
        2855 => x"cc040000",
        2856 => x"a4040000",
        2857 => x"a4040000",
        2858 => x"a4040000",
        2859 => x"a4040000",
        2860 => x"a4040000",
        2861 => x"a4040000",
        2862 => x"a4040000",
        2863 => x"a4040000",
        2864 => x"a4040000",
        2865 => x"a4040000",
        2866 => x"a4040000",
        2867 => x"a4040000",
        2868 => x"e0040000",
        2869 => x"ec040000",
        2870 => x"a8050000",
        2871 => x"90050000",
        2872 => x"a4040000",
        2873 => x"a4040000",
        2874 => x"a4040000",
        2875 => x"a4040000",
        2876 => x"a4040000",
        2877 => x"a4040000",
        2878 => x"78050000",
        2879 => x"a4040000",
        2880 => x"a4040000",
        2881 => x"a4040000",
        2882 => x"a4040000",
        2883 => x"cc040000",
        2884 => x"cc040000",
        2885 => x"00010202",
        2886 => x"03030303",
        2887 => x"04040404",
        2888 => x"04040404",
        2889 => x"05050505",
        2890 => x"05050505",
        2891 => x"05050505",
        2892 => x"05050505",
        2893 => x"06060606",
        2894 => x"06060606",
        2895 => x"06060606",
        2896 => x"06060606",
        2897 => x"06060606",
        2898 => x"06060606",
        2899 => x"06060606",
        2900 => x"06060606",
        2901 => x"07070707",
        2902 => x"07070707",
        2903 => x"07070707",
        2904 => x"07070707",
        2905 => x"07070707",
        2906 => x"07070707",
        2907 => x"07070707",
        2908 => x"07070707",
        2909 => x"07070707",
        2910 => x"07070707",
        2911 => x"07070707",
        2912 => x"07070707",
        2913 => x"07070707",
        2914 => x"07070707",
        2915 => x"07070707",
        2916 => x"07070707",
        2917 => x"08080808",
        2918 => x"08080808",
        2919 => x"08080808",
        2920 => x"08080808",
        2921 => x"08080808",
        2922 => x"08080808",
        2923 => x"08080808",
        2924 => x"08080808",
        2925 => x"08080808",
        2926 => x"08080808",
        2927 => x"08080808",
        2928 => x"08080808",
        2929 => x"08080808",
        2930 => x"08080808",
        2931 => x"08080808",
        2932 => x"08080808",
        2933 => x"08080808",
        2934 => x"08080808",
        2935 => x"08080808",
        2936 => x"08080808",
        2937 => x"08080808",
        2938 => x"08080808",
        2939 => x"08080808",
        2940 => x"08080808",
        2941 => x"08080808",
        2942 => x"08080808",
        2943 => x"08080808",
        2944 => x"08080808",
        2945 => x"08080808",
        2946 => x"08080808",
        2947 => x"08080808",
        2948 => x"08080808",
        2949 => x"0d0a4542",
        2950 => x"5245414b",
        2951 => x"21206d65",
        2952 => x"7063203d",
        2953 => x"20000000",
        2954 => x"20696e73",
        2955 => x"6e203d20",
        2956 => x"00000000",
        2957 => x"0d0a0d0a",
        2958 => x"44697370",
        2959 => x"6c617969",
        2960 => x"6e672074",
        2961 => x"68652074",
        2962 => x"696d6520",
        2963 => x"70617373",
        2964 => x"65642073",
        2965 => x"696e6365",
        2966 => x"20726573",
        2967 => x"65740d0a",
        2968 => x"0d0a0000",
        2969 => x"2530356c",
        2970 => x"643a2530",
        2971 => x"366c6420",
        2972 => x"20202530",
        2973 => x"326c643a",
        2974 => x"2530326c",
        2975 => x"643a2530",
        2976 => x"326c640d",
        2977 => x"00000000",
        2978 => x"696e7465",
        2979 => x"72727570",
        2980 => x"745f6469",
        2981 => x"72656374",
        2982 => x"00000000",
        2983 => x"54485541",
        2984 => x"53205249",
        2985 => x"53432d56",
        2986 => x"20525633",
        2987 => x"32494d20",
        2988 => x"62617265",
        2989 => x"206d6574",
        2990 => x"616c2070",
        2991 => x"726f6365",
        2992 => x"73736f72",
        2993 => x"00000000",
        2994 => x"54686520",
        2995 => x"48616775",
        2996 => x"6520556e",
        2997 => x"69766572",
        2998 => x"73697479",
        2999 => x"206f6620",
        3000 => x"4170706c",
        3001 => x"69656420",
        3002 => x"53636965",
        3003 => x"6e636573",
        3004 => x"00000000",
        3005 => x"44657061",
        3006 => x"72746d65",
        3007 => x"6e74206f",
        3008 => x"6620456c",
        3009 => x"65637472",
        3010 => x"6963616c",
        3011 => x"20456e67",
        3012 => x"696e6565",
        3013 => x"72696e67",
        3014 => x"00000000",
        3015 => x"4a2e452e",
        3016 => x"4a2e206f",
        3017 => x"70206465",
        3018 => x"6e204272",
        3019 => x"6f757700",
        3020 => x"232d302b",
        3021 => x"20000000",
        3022 => x"686c4c00",
        3023 => x"65666745",
        3024 => x"46470000",
        3025 => x"30313233",
        3026 => x"34353637",
        3027 => x"38394142",
        3028 => x"43444546",
        3029 => x"00000000",
        3030 => x"30313233",
        3031 => x"34353637",
        3032 => x"38396162",
        3033 => x"63646566",
        3034 => x"00000000",
        3035 => x"f0220000",
        3036 => x"10230000",
        3037 => x"bc220000",
        3038 => x"bc220000",
        3039 => x"bc220000",
        3040 => x"bc220000",
        3041 => x"10230000",
        3042 => x"bc220000",
        3043 => x"bc220000",
        3044 => x"bc220000",
        3045 => x"bc220000",
        3046 => x"28250000",
        3047 => x"a4230000",
        3048 => x"90240000",
        3049 => x"bc220000",
        3050 => x"bc220000",
        3051 => x"70250000",
        3052 => x"bc220000",
        3053 => x"a4230000",
        3054 => x"bc220000",
        3055 => x"bc220000",
        3056 => x"9c240000",
        3057 => x"18000020",
        3058 => x"882e0000",
        3059 => x"9c2e0000",
        3060 => x"c82e0000",
        3061 => x"f42e0000",
        3062 => x"1c2f0000",
        3063 => x"00000000",
        3064 => x"00000000",
        3065 => x"00000000",
        3066 => x"00000000",
        3067 => x"00000000",
        3068 => x"00000000",
        3069 => x"00000000",
        3070 => x"00000000",
        3071 => x"00000000",
        3072 => x"00000000",
        3073 => x"00000000",
        3074 => x"00000000",
        3075 => x"00000000",
        3076 => x"00000000",
        3077 => x"00000000",
        3078 => x"00000000",
        3079 => x"00000000",
        3080 => x"00000000",
        3081 => x"00000000",
        3082 => x"00000000",
        3083 => x"00000000",
        3084 => x"00000000",
        3085 => x"00000000",
        3086 => x"00000000",
        3087 => x"00000000",
        3088 => x"80000020",
        3089 => x"18000020",
        others => (others => '0')
    );
end package processor_common_rom;
