-- srec2vhdl table generator
-- for input file test.srec

library ieee;
use ieee.std_logic_1164.all;

library work;
use work.processor_common.all;

package processor_common_rom is
    constant rom_contents : rom_type := (
           0 => x"97110020",
           1 => x"93810180",
           2 => x"17810020",
           3 => x"130181ff",
           4 => x"97020000",
           5 => x"93828206",
           6 => x"73905230",
           7 => x"1386c187",
           8 => x"9387c188",
           9 => x"637af600",
          10 => x"3386c740",
          11 => x"93050000",
          12 => x"1385c187",
          13 => x"ef000014",
          14 => x"37050020",
          15 => x"13060500",
          16 => x"9387c187",
          17 => x"637cf600",
          18 => x"b7150000",
          19 => x"3386c740",
          20 => x"9385c56e",
          21 => x"13050500",
          22 => x"ef00800f",
          23 => x"ef000027",
          24 => x"b7050020",
          25 => x"13060000",
          26 => x"93850500",
          27 => x"13055000",
          28 => x"ef00801c",
          29 => x"ef008021",
          30 => x"6f000000",
          31 => x"b70700f0",
          32 => x"23a2a702",
          33 => x"23a4b702",
          34 => x"67800000",
          35 => x"130101ec",
          36 => x"13034112",
          37 => x"2322b112",
          38 => x"2324c112",
          39 => x"2326d112",
          40 => x"13060500",
          41 => x"93060300",
          42 => x"93050010",
          43 => x"13050101",
          44 => x"232e1110",
          45 => x"232c8110",
          46 => x"2328e112",
          47 => x"232af112",
          48 => x"232c0113",
          49 => x"232e1113",
          50 => x"23266100",
          51 => x"ef00c033",
          52 => x"13040500",
          53 => x"13050101",
          54 => x"ef008001",
          55 => x"8320c111",
          56 => x"13050400",
          57 => x"03248111",
          58 => x"13010114",
          59 => x"67800000",
          60 => x"630e0502",
          61 => x"130101ff",
          62 => x"23248100",
          63 => x"23261100",
          64 => x"13040500",
          65 => x"03450500",
          66 => x"630a0500",
          67 => x"13041400",
          68 => x"ef000002",
          69 => x"03450400",
          70 => x"e31a05fe",
          71 => x"8320c100",
          72 => x"03248100",
          73 => x"13010101",
          74 => x"67800000",
          75 => x"67800000",
          76 => x"1375f50f",
          77 => x"b70700f0",
          78 => x"23a0a702",
          79 => x"370700f0",
          80 => x"8327c702",
          81 => x"93f70701",
          82 => x"e38c07fe",
          83 => x"67800000",
          84 => x"13030500",
          85 => x"630e0600",
          86 => x"83830500",
          87 => x"23007300",
          88 => x"1306f6ff",
          89 => x"13031300",
          90 => x"93851500",
          91 => x"e31606fe",
          92 => x"67800000",
          93 => x"13030500",
          94 => x"630a0600",
          95 => x"2300b300",
          96 => x"1306f6ff",
          97 => x"13031300",
          98 => x"e31a06fe",
          99 => x"67800000",
         100 => x"630c0602",
         101 => x"13030500",
         102 => x"93061000",
         103 => x"636ab500",
         104 => x"9306f0ff",
         105 => x"1307f6ff",
         106 => x"3303e300",
         107 => x"b385e500",
         108 => x"83830500",
         109 => x"23007300",
         110 => x"1306f6ff",
         111 => x"3303d300",
         112 => x"b385d500",
         113 => x"e31606fe",
         114 => x"67800000",
         115 => x"6f000000",
         116 => x"03a7c187",
         117 => x"b7870020",
         118 => x"93870700",
         119 => x"93060040",
         120 => x"b387d740",
         121 => x"630c0700",
         122 => x"3305a700",
         123 => x"63e2a702",
         124 => x"23aea186",
         125 => x"13050700",
         126 => x"67800000",
         127 => x"93860189",
         128 => x"13870189",
         129 => x"23aed186",
         130 => x"3305a700",
         131 => x"e3f2a7fe",
         132 => x"130101ff",
         133 => x"23261100",
         134 => x"ef104038",
         135 => x"8320c100",
         136 => x"9307c000",
         137 => x"2320f500",
         138 => x"1307f0ff",
         139 => x"13050700",
         140 => x"13010101",
         141 => x"67800000",
         142 => x"b7676c6c",
         143 => x"130101fe",
         144 => x"93878754",
         145 => x"2324f100",
         146 => x"93050000",
         147 => x"9307f006",
         148 => x"1305101b",
         149 => x"232e1100",
         150 => x"2316f100",
         151 => x"eff01fe2",
         152 => x"93068100",
         153 => x"37150000",
         154 => x"1307f00f",
         155 => x"13063000",
         156 => x"93850600",
         157 => x"13050564",
         158 => x"eff05fe1",
         159 => x"8320c101",
         160 => x"13050000",
         161 => x"13010102",
         162 => x"67800000",
         163 => x"130101ff",
         164 => x"23248100",
         165 => x"23261100",
         166 => x"93070000",
         167 => x"13040500",
         168 => x"63880700",
         169 => x"93050000",
         170 => x"97000000",
         171 => x"e7000000",
         172 => x"b7170000",
         173 => x"03a5876e",
         174 => x"83278502",
         175 => x"63840700",
         176 => x"e7800700",
         177 => x"13050400",
         178 => x"eff05ff0",
         179 => x"130101ff",
         180 => x"23248100",
         181 => x"23229100",
         182 => x"37140000",
         183 => x"b7140000",
         184 => x"9387c46e",
         185 => x"1304c46e",
         186 => x"3304f440",
         187 => x"23202101",
         188 => x"23261100",
         189 => x"13542440",
         190 => x"9384c46e",
         191 => x"13090000",
         192 => x"63108904",
         193 => x"b7140000",
         194 => x"37140000",
         195 => x"9387c46e",
         196 => x"1304c46e",
         197 => x"3304f440",
         198 => x"13542440",
         199 => x"9384c46e",
         200 => x"13090000",
         201 => x"63188902",
         202 => x"8320c100",
         203 => x"03248100",
         204 => x"83244100",
         205 => x"03290100",
         206 => x"13010101",
         207 => x"67800000",
         208 => x"83a70400",
         209 => x"13091900",
         210 => x"93844400",
         211 => x"e7800700",
         212 => x"6ff01ffb",
         213 => x"83a70400",
         214 => x"13091900",
         215 => x"93844400",
         216 => x"e7800700",
         217 => x"6ff01ffc",
         218 => x"130101f8",
         219 => x"232c8106",
         220 => x"232a9106",
         221 => x"232e1106",
         222 => x"23282107",
         223 => x"93040500",
         224 => x"13040600",
         225 => x"63540602",
         226 => x"9307b008",
         227 => x"2320f500",
         228 => x"1305f0ff",
         229 => x"8320c107",
         230 => x"03248107",
         231 => x"83244107",
         232 => x"03290107",
         233 => x"13010108",
         234 => x"67800000",
         235 => x"93078020",
         236 => x"231af100",
         237 => x"2324b100",
         238 => x"232cb100",
         239 => x"13860600",
         240 => x"93070000",
         241 => x"93060700",
         242 => x"63040400",
         243 => x"9307f4ff",
         244 => x"1309f0ff",
         245 => x"93058100",
         246 => x"13850400",
         247 => x"2328f100",
         248 => x"232ef100",
         249 => x"231b2101",
         250 => x"ef000036",
         251 => x"63562501",
         252 => x"9307b008",
         253 => x"23a0f400",
         254 => x"e30e04f8",
         255 => x"83278100",
         256 => x"23800700",
         257 => x"6ff01ff9",
         258 => x"13870600",
         259 => x"93060600",
         260 => x"13860500",
         261 => x"93050500",
         262 => x"03a58187",
         263 => x"6ff0dff4",
         264 => x"130101fe",
         265 => x"23282101",
         266 => x"03a98500",
         267 => x"232c8100",
         268 => x"23263101",
         269 => x"23225101",
         270 => x"23206101",
         271 => x"232e1100",
         272 => x"232a9100",
         273 => x"23244101",
         274 => x"83aa0500",
         275 => x"13840500",
         276 => x"130b0600",
         277 => x"93890600",
         278 => x"63ec2609",
         279 => x"8397c500",
         280 => x"13f70748",
         281 => x"63040708",
         282 => x"03274401",
         283 => x"93043000",
         284 => x"83a50501",
         285 => x"b384e402",
         286 => x"13072000",
         287 => x"b38aba40",
         288 => x"130a0500",
         289 => x"b3c4e402",
         290 => x"13871600",
         291 => x"33075701",
         292 => x"63f4e400",
         293 => x"93040700",
         294 => x"93f70740",
         295 => x"6386070a",
         296 => x"93850400",
         297 => x"13050a00",
         298 => x"ef00104c",
         299 => x"13090500",
         300 => x"630c050a",
         301 => x"83250401",
         302 => x"13860a00",
         303 => x"eff05fc9",
         304 => x"8357c400",
         305 => x"93f7f7b7",
         306 => x"93e70708",
         307 => x"2316f400",
         308 => x"23282401",
         309 => x"232a9400",
         310 => x"33095901",
         311 => x"b3845441",
         312 => x"23202401",
         313 => x"23249400",
         314 => x"13890900",
         315 => x"63f42901",
         316 => x"13890900",
         317 => x"03250400",
         318 => x"13060900",
         319 => x"93050b00",
         320 => x"eff01fc9",
         321 => x"83278400",
         322 => x"13050000",
         323 => x"b3872741",
         324 => x"2324f400",
         325 => x"83270400",
         326 => x"b3872701",
         327 => x"2320f400",
         328 => x"8320c101",
         329 => x"03248101",
         330 => x"83244101",
         331 => x"03290101",
         332 => x"8329c100",
         333 => x"032a8100",
         334 => x"832a4100",
         335 => x"032b0100",
         336 => x"13010102",
         337 => x"67800000",
         338 => x"13860400",
         339 => x"13050a00",
         340 => x"ef001056",
         341 => x"13090500",
         342 => x"e31c05f6",
         343 => x"83250401",
         344 => x"13050a00",
         345 => x"ef00d030",
         346 => x"9307c000",
         347 => x"2320fa00",
         348 => x"8357c400",
         349 => x"1305f0ff",
         350 => x"93e70704",
         351 => x"2316f400",
         352 => x"6ff01ffa",
         353 => x"83278600",
         354 => x"130101fd",
         355 => x"232e3101",
         356 => x"23286101",
         357 => x"23261102",
         358 => x"23248102",
         359 => x"23229102",
         360 => x"23202103",
         361 => x"232c4101",
         362 => x"232a5101",
         363 => x"23267101",
         364 => x"23248101",
         365 => x"23229101",
         366 => x"2320a101",
         367 => x"032b0600",
         368 => x"93090600",
         369 => x"63940712",
         370 => x"13050000",
         371 => x"8320c102",
         372 => x"03248102",
         373 => x"23a20900",
         374 => x"83244102",
         375 => x"03290102",
         376 => x"8329c101",
         377 => x"032a8101",
         378 => x"832a4101",
         379 => x"032b0101",
         380 => x"832bc100",
         381 => x"032c8100",
         382 => x"832c4100",
         383 => x"032d0100",
         384 => x"13010103",
         385 => x"67800000",
         386 => x"832b0b00",
         387 => x"032d4b00",
         388 => x"130b8b00",
         389 => x"03298400",
         390 => x"832a0400",
         391 => x"e3060dfe",
         392 => x"63642d09",
         393 => x"8317c400",
         394 => x"13f70748",
         395 => x"630e0706",
         396 => x"83244401",
         397 => x"83250401",
         398 => x"b3049c02",
         399 => x"b38aba40",
         400 => x"13871a00",
         401 => x"3307a701",
         402 => x"b3c49403",
         403 => x"63f4e400",
         404 => x"93040700",
         405 => x"93f70740",
         406 => x"6388070a",
         407 => x"93850400",
         408 => x"13050a00",
         409 => x"ef005030",
         410 => x"13090500",
         411 => x"630e050a",
         412 => x"83250401",
         413 => x"13860a00",
         414 => x"eff09fad",
         415 => x"8357c400",
         416 => x"93f7f7b7",
         417 => x"93e70708",
         418 => x"2316f400",
         419 => x"23282401",
         420 => x"232a9400",
         421 => x"33095901",
         422 => x"b3845441",
         423 => x"23202401",
         424 => x"23249400",
         425 => x"13090d00",
         426 => x"63742d01",
         427 => x"13090d00",
         428 => x"03250400",
         429 => x"13060900",
         430 => x"93850b00",
         431 => x"eff05fad",
         432 => x"83278400",
         433 => x"b3872741",
         434 => x"2324f400",
         435 => x"83270400",
         436 => x"b3872701",
         437 => x"2320f400",
         438 => x"83a78900",
         439 => x"b387a741",
         440 => x"23a4f900",
         441 => x"e39207f2",
         442 => x"6ff01fee",
         443 => x"130a0500",
         444 => x"13840500",
         445 => x"930b0000",
         446 => x"130d0000",
         447 => x"130c3000",
         448 => x"930c2000",
         449 => x"6ff01ff1",
         450 => x"13860400",
         451 => x"13050a00",
         452 => x"ef00103a",
         453 => x"13090500",
         454 => x"e31a05f6",
         455 => x"83250401",
         456 => x"13050a00",
         457 => x"ef00d014",
         458 => x"9307c000",
         459 => x"2320fa00",
         460 => x"8357c400",
         461 => x"1305f0ff",
         462 => x"93e70704",
         463 => x"2316f400",
         464 => x"23a40900",
         465 => x"6ff09fe8",
         466 => x"83d7c500",
         467 => x"130101f5",
         468 => x"2324810a",
         469 => x"2322910a",
         470 => x"2320210b",
         471 => x"232c4109",
         472 => x"2326110a",
         473 => x"232e3109",
         474 => x"232a5109",
         475 => x"23286109",
         476 => x"23267109",
         477 => x"23248109",
         478 => x"23229109",
         479 => x"2320a109",
         480 => x"232eb107",
         481 => x"93f70708",
         482 => x"130a0500",
         483 => x"13890500",
         484 => x"93040600",
         485 => x"13840600",
         486 => x"63880706",
         487 => x"83a70501",
         488 => x"63940706",
         489 => x"93050004",
         490 => x"ef00101c",
         491 => x"2320a900",
         492 => x"2328a900",
         493 => x"63160504",
         494 => x"9307c000",
         495 => x"2320fa00",
         496 => x"1305f0ff",
         497 => x"8320c10a",
         498 => x"0324810a",
         499 => x"8324410a",
         500 => x"0329010a",
         501 => x"8329c109",
         502 => x"032a8109",
         503 => x"832a4109",
         504 => x"032b0109",
         505 => x"832bc108",
         506 => x"032c8108",
         507 => x"832c4108",
         508 => x"032d0108",
         509 => x"832dc107",
         510 => x"1301010b",
         511 => x"67800000",
         512 => x"93070004",
         513 => x"232af900",
         514 => x"93070002",
         515 => x"a304f102",
         516 => x"93070003",
         517 => x"23220102",
         518 => x"2305f102",
         519 => x"23268100",
         520 => x"930c5002",
         521 => x"371b0000",
         522 => x"b71b0000",
         523 => x"371d0000",
         524 => x"930a0000",
         525 => x"13840400",
         526 => x"83470400",
         527 => x"63840700",
         528 => x"639c970d",
         529 => x"b30d9440",
         530 => x"63069402",
         531 => x"93860d00",
         532 => x"13860400",
         533 => x"93050900",
         534 => x"13050a00",
         535 => x"eff05fbc",
         536 => x"9307f0ff",
         537 => x"6304f524",
         538 => x"83274102",
         539 => x"b387b701",
         540 => x"2322f102",
         541 => x"83470400",
         542 => x"638a0722",
         543 => x"9307f0ff",
         544 => x"93041400",
         545 => x"23280100",
         546 => x"232e0100",
         547 => x"232af100",
         548 => x"232c0100",
         549 => x"a3090104",
         550 => x"23240106",
         551 => x"930d1000",
         552 => x"83c50400",
         553 => x"13065000",
         554 => x"13054b65",
         555 => x"ef00007a",
         556 => x"83270101",
         557 => x"13841400",
         558 => x"63140506",
         559 => x"13f70701",
         560 => x"63060700",
         561 => x"13070002",
         562 => x"a309e104",
         563 => x"13f78700",
         564 => x"63060700",
         565 => x"1307b002",
         566 => x"a309e104",
         567 => x"83c60400",
         568 => x"1307a002",
         569 => x"638ce604",
         570 => x"8327c101",
         571 => x"13840400",
         572 => x"93060000",
         573 => x"13069000",
         574 => x"1305a000",
         575 => x"03470400",
         576 => x"93051400",
         577 => x"130707fd",
         578 => x"637ee608",
         579 => x"63840604",
         580 => x"232ef100",
         581 => x"6f000004",
         582 => x"13041400",
         583 => x"6ff0dff1",
         584 => x"13074b65",
         585 => x"3305e540",
         586 => x"3395ad00",
         587 => x"b3e7a700",
         588 => x"2328f100",
         589 => x"93040400",
         590 => x"6ff09ff6",
         591 => x"0327c100",
         592 => x"93064700",
         593 => x"03270700",
         594 => x"2326d100",
         595 => x"63420704",
         596 => x"232ee100",
         597 => x"03470400",
         598 => x"9307e002",
         599 => x"6314f708",
         600 => x"03471400",
         601 => x"9307a002",
         602 => x"6318f704",
         603 => x"8327c100",
         604 => x"13042400",
         605 => x"13874700",
         606 => x"83a70700",
         607 => x"2326e100",
         608 => x"63d40700",
         609 => x"9307f0ff",
         610 => x"232af100",
         611 => x"6f008005",
         612 => x"3307e040",
         613 => x"93e72700",
         614 => x"232ee100",
         615 => x"2328f100",
         616 => x"6ff05ffb",
         617 => x"b387a702",
         618 => x"13840500",
         619 => x"93061000",
         620 => x"b387e700",
         621 => x"6ff09ff4",
         622 => x"13041400",
         623 => x"232a0100",
         624 => x"93060000",
         625 => x"93070000",
         626 => x"13069000",
         627 => x"1305a000",
         628 => x"03470400",
         629 => x"93051400",
         630 => x"130707fd",
         631 => x"6372e608",
         632 => x"e39406fa",
         633 => x"83450400",
         634 => x"13063000",
         635 => x"1385cb65",
         636 => x"ef00c065",
         637 => x"63020502",
         638 => x"9387cb65",
         639 => x"3305f540",
         640 => x"83270101",
         641 => x"13070004",
         642 => x"3317a700",
         643 => x"b3e7e700",
         644 => x"13041400",
         645 => x"2328f100",
         646 => x"83450400",
         647 => x"13066000",
         648 => x"13050d66",
         649 => x"93041400",
         650 => x"2304b102",
         651 => x"ef000062",
         652 => x"63080508",
         653 => x"63980a04",
         654 => x"03270101",
         655 => x"8327c100",
         656 => x"13770710",
         657 => x"63080702",
         658 => x"93874700",
         659 => x"2326f100",
         660 => x"83274102",
         661 => x"b3873701",
         662 => x"2322f102",
         663 => x"6ff09fdd",
         664 => x"b387a702",
         665 => x"13840500",
         666 => x"93061000",
         667 => x"b387e700",
         668 => x"6ff01ff6",
         669 => x"93877700",
         670 => x"93f787ff",
         671 => x"93878700",
         672 => x"6ff0dffc",
         673 => x"1307c100",
         674 => x"93060042",
         675 => x"13060900",
         676 => x"93050101",
         677 => x"13050a00",
         678 => x"97000000",
         679 => x"e7000000",
         680 => x"9307f0ff",
         681 => x"93090500",
         682 => x"e314f5fa",
         683 => x"8357c900",
         684 => x"93f70704",
         685 => x"e39607d0",
         686 => x"03254102",
         687 => x"6ff09fd0",
         688 => x"1307c100",
         689 => x"93060042",
         690 => x"13060900",
         691 => x"93050101",
         692 => x"13050a00",
         693 => x"ef00801b",
         694 => x"6ff09ffc",
         695 => x"130101fd",
         696 => x"232a5101",
         697 => x"83a70501",
         698 => x"930a0700",
         699 => x"03a78500",
         700 => x"23248102",
         701 => x"23202103",
         702 => x"232e3101",
         703 => x"232c4101",
         704 => x"23261102",
         705 => x"23229102",
         706 => x"23286101",
         707 => x"23267101",
         708 => x"93090500",
         709 => x"13840500",
         710 => x"13090600",
         711 => x"138a0600",
         712 => x"63d4e700",
         713 => x"93070700",
         714 => x"2320f900",
         715 => x"03473404",
         716 => x"63060700",
         717 => x"93871700",
         718 => x"2320f900",
         719 => x"83270400",
         720 => x"93f70702",
         721 => x"63880700",
         722 => x"83270900",
         723 => x"93872700",
         724 => x"2320f900",
         725 => x"83240400",
         726 => x"93f46400",
         727 => x"639e0400",
         728 => x"130b9401",
         729 => x"930bf0ff",
         730 => x"8327c400",
         731 => x"03270900",
         732 => x"b387e740",
         733 => x"63c2f408",
         734 => x"83473404",
         735 => x"b336f000",
         736 => x"83270400",
         737 => x"93f70702",
         738 => x"6390070c",
         739 => x"13063404",
         740 => x"93050a00",
         741 => x"13850900",
         742 => x"e7800a00",
         743 => x"9307f0ff",
         744 => x"6308f506",
         745 => x"83270400",
         746 => x"13074000",
         747 => x"93040000",
         748 => x"93f76700",
         749 => x"639ce700",
         750 => x"8324c400",
         751 => x"83270900",
         752 => x"b384f440",
         753 => x"63d40400",
         754 => x"93040000",
         755 => x"83278400",
         756 => x"03270401",
         757 => x"6356f700",
         758 => x"b387e740",
         759 => x"b384f400",
         760 => x"13090000",
         761 => x"1304a401",
         762 => x"130bf0ff",
         763 => x"63902409",
         764 => x"13050000",
         765 => x"6f000002",
         766 => x"93061000",
         767 => x"13060b00",
         768 => x"93050a00",
         769 => x"13850900",
         770 => x"e7800a00",
         771 => x"631a7503",
         772 => x"1305f0ff",
         773 => x"8320c102",
         774 => x"03248102",
         775 => x"83244102",
         776 => x"03290102",
         777 => x"8329c101",
         778 => x"032a8101",
         779 => x"832a4101",
         780 => x"032b0101",
         781 => x"832bc100",
         782 => x"13010103",
         783 => x"67800000",
         784 => x"93841400",
         785 => x"6ff05ff2",
         786 => x"3307d400",
         787 => x"13060003",
         788 => x"a301c704",
         789 => x"03475404",
         790 => x"93871600",
         791 => x"b307f400",
         792 => x"93862600",
         793 => x"a381e704",
         794 => x"6ff05ff2",
         795 => x"93061000",
         796 => x"13060400",
         797 => x"93050a00",
         798 => x"13850900",
         799 => x"e7800a00",
         800 => x"e30865f9",
         801 => x"13091900",
         802 => x"6ff05ff6",
         803 => x"130101fd",
         804 => x"23248102",
         805 => x"23229102",
         806 => x"23202103",
         807 => x"232e3101",
         808 => x"23261102",
         809 => x"232c4101",
         810 => x"232a5101",
         811 => x"23286101",
         812 => x"83c88501",
         813 => x"93078007",
         814 => x"93040500",
         815 => x"13840500",
         816 => x"13090600",
         817 => x"93890600",
         818 => x"63ee1701",
         819 => x"93072006",
         820 => x"93863504",
         821 => x"63ee1701",
         822 => x"638a082a",
         823 => x"93078005",
         824 => x"638af820",
         825 => x"930a2404",
         826 => x"23011405",
         827 => x"6f004004",
         828 => x"9387d8f9",
         829 => x"93f7f70f",
         830 => x"13065001",
         831 => x"e364f6fe",
         832 => x"37160000",
         833 => x"93972700",
         834 => x"13060669",
         835 => x"b387c700",
         836 => x"83a70700",
         837 => x"67800700",
         838 => x"83270700",
         839 => x"938a2504",
         840 => x"93864700",
         841 => x"83a70700",
         842 => x"2320d700",
         843 => x"2381f504",
         844 => x"93071000",
         845 => x"6f004029",
         846 => x"03a60500",
         847 => x"83270700",
         848 => x"13750608",
         849 => x"93854700",
         850 => x"630e0504",
         851 => x"83a70700",
         852 => x"2320b700",
         853 => x"37170000",
         854 => x"83254400",
         855 => x"13088766",
         856 => x"63d2071e",
         857 => x"1307d002",
         858 => x"a301e404",
         859 => x"2324b400",
         860 => x"63d80504",
         861 => x"b307f040",
         862 => x"1307a000",
         863 => x"938a0600",
         864 => x"33f6e702",
         865 => x"938afaff",
         866 => x"3306c800",
         867 => x"03460600",
         868 => x"2380ca00",
         869 => x"13860700",
         870 => x"b3d7e702",
         871 => x"e372e6fe",
         872 => x"6f008009",
         873 => x"83a70700",
         874 => x"13750604",
         875 => x"2320b700",
         876 => x"e30205fa",
         877 => x"93970701",
         878 => x"93d70741",
         879 => x"6ff09ff9",
         880 => x"1376b6ff",
         881 => x"2320c400",
         882 => x"6ff0dffa",
         883 => x"03a60500",
         884 => x"83270700",
         885 => x"13750608",
         886 => x"93854700",
         887 => x"63080500",
         888 => x"2320b700",
         889 => x"83a70700",
         890 => x"6f004001",
         891 => x"13760604",
         892 => x"2320b700",
         893 => x"e30806fe",
         894 => x"83d70700",
         895 => x"37180000",
         896 => x"1307f006",
         897 => x"13088866",
         898 => x"639ae812",
         899 => x"13078000",
         900 => x"a3010404",
         901 => x"03264400",
         902 => x"2324c400",
         903 => x"e34006f6",
         904 => x"83250400",
         905 => x"93f5b5ff",
         906 => x"2320b400",
         907 => x"e39807f4",
         908 => x"938a0600",
         909 => x"e31406f4",
         910 => x"93078000",
         911 => x"6314f702",
         912 => x"83270400",
         913 => x"93f71700",
         914 => x"638e0700",
         915 => x"03274400",
         916 => x"83270401",
         917 => x"63c8e700",
         918 => x"93070003",
         919 => x"a38ffafe",
         920 => x"938afaff",
         921 => x"b3865641",
         922 => x"2328d400",
         923 => x"13870900",
         924 => x"93060900",
         925 => x"1306c100",
         926 => x"93050400",
         927 => x"13850400",
         928 => x"eff0dfc5",
         929 => x"130af0ff",
         930 => x"63164515",
         931 => x"1305f0ff",
         932 => x"8320c102",
         933 => x"03248102",
         934 => x"83244102",
         935 => x"03290102",
         936 => x"8329c101",
         937 => x"032a8101",
         938 => x"832a4101",
         939 => x"032b0101",
         940 => x"13010103",
         941 => x"67800000",
         942 => x"83a70500",
         943 => x"93e70702",
         944 => x"23a0f500",
         945 => x"37180000",
         946 => x"93088007",
         947 => x"1308c867",
         948 => x"03260400",
         949 => x"a3021405",
         950 => x"83270700",
         951 => x"13750608",
         952 => x"93854700",
         953 => x"630e0500",
         954 => x"2320b700",
         955 => x"83a70700",
         956 => x"6f000002",
         957 => x"37180000",
         958 => x"13088866",
         959 => x"6ff05ffd",
         960 => x"13750604",
         961 => x"2320b700",
         962 => x"e30205fe",
         963 => x"83d70700",
         964 => x"13771600",
         965 => x"63060700",
         966 => x"13660602",
         967 => x"2320c400",
         968 => x"63860700",
         969 => x"13070001",
         970 => x"6ff09fee",
         971 => x"03270400",
         972 => x"1377f7fd",
         973 => x"2320e400",
         974 => x"6ff0dffe",
         975 => x"1307a000",
         976 => x"6ff01fed",
         977 => x"13088766",
         978 => x"1307a000",
         979 => x"6ff09fec",
         980 => x"03a60500",
         981 => x"83270700",
         982 => x"83a54501",
         983 => x"13780608",
         984 => x"13854700",
         985 => x"630a0800",
         986 => x"2320a700",
         987 => x"83a70700",
         988 => x"23a0b700",
         989 => x"6f008001",
         990 => x"2320a700",
         991 => x"13760604",
         992 => x"83a70700",
         993 => x"e30606fe",
         994 => x"2390b700",
         995 => x"23280400",
         996 => x"938a0600",
         997 => x"6ff09fed",
         998 => x"83270700",
         999 => x"03a64500",
        1000 => x"93050000",
        1001 => x"93864700",
        1002 => x"2320d700",
        1003 => x"83aa0700",
        1004 => x"13850a00",
        1005 => x"ef008009",
        1006 => x"63060500",
        1007 => x"33055541",
        1008 => x"2322a400",
        1009 => x"83274400",
        1010 => x"2328f400",
        1011 => x"a3010404",
        1012 => x"6ff0dfe9",
        1013 => x"83260401",
        1014 => x"13860a00",
        1015 => x"93050900",
        1016 => x"13850400",
        1017 => x"e7800900",
        1018 => x"e30245eb",
        1019 => x"83270400",
        1020 => x"93f72700",
        1021 => x"63940704",
        1022 => x"8327c100",
        1023 => x"0325c400",
        1024 => x"e358f5e8",
        1025 => x"13850700",
        1026 => x"6ff09fe8",
        1027 => x"93061000",
        1028 => x"13860a00",
        1029 => x"93050900",
        1030 => x"13850400",
        1031 => x"e7800900",
        1032 => x"e30665e7",
        1033 => x"130a1a00",
        1034 => x"8327c400",
        1035 => x"0327c100",
        1036 => x"b387e740",
        1037 => x"e34cfafc",
        1038 => x"6ff01ffc",
        1039 => x"130a0000",
        1040 => x"930a9401",
        1041 => x"130bf0ff",
        1042 => x"6ff01ffe",
        1043 => x"93f5f50f",
        1044 => x"3306c500",
        1045 => x"6316c500",
        1046 => x"13050000",
        1047 => x"67800000",
        1048 => x"83470500",
        1049 => x"e38cb7fe",
        1050 => x"13051500",
        1051 => x"6ff09ffe",
        1052 => x"638a050e",
        1053 => x"83a7c5ff",
        1054 => x"130101fe",
        1055 => x"232c8100",
        1056 => x"232e1100",
        1057 => x"1384c5ff",
        1058 => x"63d40700",
        1059 => x"3304f400",
        1060 => x"2326a100",
        1061 => x"ef008033",
        1062 => x"83a74188",
        1063 => x"0325c100",
        1064 => x"639e0700",
        1065 => x"23220400",
        1066 => x"23a28188",
        1067 => x"03248101",
        1068 => x"8320c101",
        1069 => x"13010102",
        1070 => x"6f008031",
        1071 => x"6374f402",
        1072 => x"03260400",
        1073 => x"b306c400",
        1074 => x"639ad700",
        1075 => x"83a60700",
        1076 => x"83a74700",
        1077 => x"b386c600",
        1078 => x"2320d400",
        1079 => x"2322f400",
        1080 => x"6ff09ffc",
        1081 => x"13870700",
        1082 => x"83a74700",
        1083 => x"63840700",
        1084 => x"e37af4fe",
        1085 => x"83260700",
        1086 => x"3306d700",
        1087 => x"63188602",
        1088 => x"03260400",
        1089 => x"b386c600",
        1090 => x"2320d700",
        1091 => x"3306d700",
        1092 => x"e39ec7f8",
        1093 => x"03a60700",
        1094 => x"83a74700",
        1095 => x"b306d600",
        1096 => x"2320d700",
        1097 => x"2322f700",
        1098 => x"6ff05ff8",
        1099 => x"6378c400",
        1100 => x"9307c000",
        1101 => x"2320f500",
        1102 => x"6ff05ff7",
        1103 => x"03260400",
        1104 => x"b306c400",
        1105 => x"639ad700",
        1106 => x"83a60700",
        1107 => x"83a74700",
        1108 => x"b386c600",
        1109 => x"2320d400",
        1110 => x"2322f400",
        1111 => x"23228700",
        1112 => x"6ff0dff4",
        1113 => x"67800000",
        1114 => x"130101fe",
        1115 => x"232a9100",
        1116 => x"93843500",
        1117 => x"93f4c4ff",
        1118 => x"23282101",
        1119 => x"232e1100",
        1120 => x"232c8100",
        1121 => x"23263101",
        1122 => x"93848400",
        1123 => x"9307c000",
        1124 => x"13090500",
        1125 => x"63f0f406",
        1126 => x"9304c000",
        1127 => x"63eeb404",
        1128 => x"13050900",
        1129 => x"ef008022",
        1130 => x"03a74188",
        1131 => x"13040700",
        1132 => x"63180406",
        1133 => x"83a70188",
        1134 => x"639a0700",
        1135 => x"93050000",
        1136 => x"13050900",
        1137 => x"ef00001c",
        1138 => x"23a0a188",
        1139 => x"93850400",
        1140 => x"13050900",
        1141 => x"ef00001b",
        1142 => x"9309f0ff",
        1143 => x"631a350b",
        1144 => x"9307c000",
        1145 => x"2320f900",
        1146 => x"13050900",
        1147 => x"ef00401e",
        1148 => x"6f000001",
        1149 => x"e3d404fa",
        1150 => x"9307c000",
        1151 => x"2320f900",
        1152 => x"13050000",
        1153 => x"8320c101",
        1154 => x"03248101",
        1155 => x"83244101",
        1156 => x"03290101",
        1157 => x"8329c100",
        1158 => x"13010102",
        1159 => x"67800000",
        1160 => x"83270400",
        1161 => x"b3879740",
        1162 => x"63ce0704",
        1163 => x"1306b000",
        1164 => x"637af600",
        1165 => x"2320f400",
        1166 => x"3304f400",
        1167 => x"23209400",
        1168 => x"6f000001",
        1169 => x"83274400",
        1170 => x"631a8702",
        1171 => x"23a2f188",
        1172 => x"13050900",
        1173 => x"ef00c017",
        1174 => x"1305b400",
        1175 => x"93074400",
        1176 => x"137585ff",
        1177 => x"3307f540",
        1178 => x"e30ef5f8",
        1179 => x"3304e400",
        1180 => x"b387a740",
        1181 => x"2320f400",
        1182 => x"6ff0dff8",
        1183 => x"2322f700",
        1184 => x"6ff01ffd",
        1185 => x"13070400",
        1186 => x"03244400",
        1187 => x"6ff05ff2",
        1188 => x"13043500",
        1189 => x"1374c4ff",
        1190 => x"e30285fa",
        1191 => x"b305a440",
        1192 => x"13050900",
        1193 => x"ef00000e",
        1194 => x"e31a35f9",
        1195 => x"6ff05ff3",
        1196 => x"130101fe",
        1197 => x"232c8100",
        1198 => x"232e1100",
        1199 => x"232a9100",
        1200 => x"23282101",
        1201 => x"23263101",
        1202 => x"23244101",
        1203 => x"13040600",
        1204 => x"63940502",
        1205 => x"03248101",
        1206 => x"8320c101",
        1207 => x"83244101",
        1208 => x"03290101",
        1209 => x"8329c100",
        1210 => x"032a8100",
        1211 => x"93050600",
        1212 => x"13010102",
        1213 => x"6ff05fe7",
        1214 => x"63180602",
        1215 => x"eff05fd7",
        1216 => x"93040000",
        1217 => x"8320c101",
        1218 => x"03248101",
        1219 => x"03290101",
        1220 => x"8329c100",
        1221 => x"032a8100",
        1222 => x"13850400",
        1223 => x"83244101",
        1224 => x"13010102",
        1225 => x"67800000",
        1226 => x"130a0500",
        1227 => x"93840500",
        1228 => x"ef00400a",
        1229 => x"13090500",
        1230 => x"63668500",
        1231 => x"93571500",
        1232 => x"e3e287fc",
        1233 => x"93050400",
        1234 => x"13050a00",
        1235 => x"eff0dfe1",
        1236 => x"93090500",
        1237 => x"e30605fa",
        1238 => x"13060400",
        1239 => x"63748900",
        1240 => x"13060900",
        1241 => x"93850400",
        1242 => x"13850900",
        1243 => x"efe05fde",
        1244 => x"93850400",
        1245 => x"13050a00",
        1246 => x"eff09fcf",
        1247 => x"93840900",
        1248 => x"6ff05ff8",
        1249 => x"130101ff",
        1250 => x"23248100",
        1251 => x"23229100",
        1252 => x"13040500",
        1253 => x"13850500",
        1254 => x"23261100",
        1255 => x"23a40188",
        1256 => x"efe01fe3",
        1257 => x"9307f0ff",
        1258 => x"6318f500",
        1259 => x"83a78188",
        1260 => x"63840700",
        1261 => x"2320f400",
        1262 => x"8320c100",
        1263 => x"03248100",
        1264 => x"83244100",
        1265 => x"13010101",
        1266 => x"67800000",
        1267 => x"67800000",
        1268 => x"67800000",
        1269 => x"83a7c5ff",
        1270 => x"1385c7ff",
        1271 => x"63d80700",
        1272 => x"b385a500",
        1273 => x"83a70500",
        1274 => x"3305f500",
        1275 => x"67800000",
        1276 => x"130101ff",
        1277 => x"23248100",
        1278 => x"13840500",
        1279 => x"83a50500",
        1280 => x"23229100",
        1281 => x"23261100",
        1282 => x"93040500",
        1283 => x"63840500",
        1284 => x"eff01ffe",
        1285 => x"93050400",
        1286 => x"03248100",
        1287 => x"8320c100",
        1288 => x"13850400",
        1289 => x"83244100",
        1290 => x"13010101",
        1291 => x"6ff05fc4",
        1292 => x"83a78187",
        1293 => x"6382a716",
        1294 => x"83274502",
        1295 => x"130101fe",
        1296 => x"232c8100",
        1297 => x"232e1100",
        1298 => x"232a9100",
        1299 => x"23282101",
        1300 => x"23263101",
        1301 => x"13040500",
        1302 => x"638a0704",
        1303 => x"83a7c700",
        1304 => x"638c0702",
        1305 => x"93040000",
        1306 => x"13090008",
        1307 => x"83274402",
        1308 => x"83a7c700",
        1309 => x"b3879700",
        1310 => x"83a50700",
        1311 => x"6396050e",
        1312 => x"93844400",
        1313 => x"e39424ff",
        1314 => x"83274402",
        1315 => x"13050400",
        1316 => x"83a5c700",
        1317 => x"eff0dfbd",
        1318 => x"83274402",
        1319 => x"83a50700",
        1320 => x"63860500",
        1321 => x"13050400",
        1322 => x"eff09fbc",
        1323 => x"83254401",
        1324 => x"63860500",
        1325 => x"13050400",
        1326 => x"eff09fbb",
        1327 => x"83254402",
        1328 => x"63860500",
        1329 => x"13050400",
        1330 => x"eff09fba",
        1331 => x"83258403",
        1332 => x"63860500",
        1333 => x"13050400",
        1334 => x"eff09fb9",
        1335 => x"8325c403",
        1336 => x"63860500",
        1337 => x"13050400",
        1338 => x"eff09fb8",
        1339 => x"83250404",
        1340 => x"63860500",
        1341 => x"13050400",
        1342 => x"eff09fb7",
        1343 => x"8325c405",
        1344 => x"63860500",
        1345 => x"13050400",
        1346 => x"eff09fb6",
        1347 => x"83258405",
        1348 => x"63860500",
        1349 => x"13050400",
        1350 => x"eff09fb5",
        1351 => x"83254403",
        1352 => x"63860500",
        1353 => x"13050400",
        1354 => x"eff09fb4",
        1355 => x"83278401",
        1356 => x"63860704",
        1357 => x"83278402",
        1358 => x"13050400",
        1359 => x"e7800700",
        1360 => x"83258404",
        1361 => x"638c0502",
        1362 => x"13050400",
        1363 => x"03248101",
        1364 => x"8320c101",
        1365 => x"83244101",
        1366 => x"03290101",
        1367 => x"8329c100",
        1368 => x"13010102",
        1369 => x"6ff0dfe8",
        1370 => x"83a90500",
        1371 => x"13050400",
        1372 => x"eff01fb0",
        1373 => x"93850900",
        1374 => x"6ff05ff0",
        1375 => x"8320c101",
        1376 => x"03248101",
        1377 => x"83244101",
        1378 => x"03290101",
        1379 => x"8329c100",
        1380 => x"13010102",
        1381 => x"67800000",
        1382 => x"67800000",
        1383 => x"03a58187",
        1384 => x"67800000",
        1385 => x"74657374",
        1386 => x"00000000",
        1387 => x"54485541",
        1388 => x"53205249",
        1389 => x"53432d56",
        1390 => x"20525633",
        1391 => x"32494d20",
        1392 => x"62617265",
        1393 => x"206d6574",
        1394 => x"616c2070",
        1395 => x"726f6365",
        1396 => x"73736f72",
        1397 => x"00000000",
        1398 => x"54686520",
        1399 => x"48616775",
        1400 => x"6520556e",
        1401 => x"69766572",
        1402 => x"73697479",
        1403 => x"206f6620",
        1404 => x"4170706c",
        1405 => x"69656420",
        1406 => x"53636965",
        1407 => x"6e636573",
        1408 => x"00000000",
        1409 => x"44657061",
        1410 => x"72746d65",
        1411 => x"6e74206f",
        1412 => x"6620456c",
        1413 => x"65637472",
        1414 => x"6963616c",
        1415 => x"20456e67",
        1416 => x"696e6565",
        1417 => x"72696e67",
        1418 => x"00000000",
        1419 => x"4a2e452e",
        1420 => x"4a2e206f",
        1421 => x"70206465",
        1422 => x"6e204272",
        1423 => x"6f757700",
        1424 => x"25732c20",
        1425 => x"25642c20",
        1426 => x"25702c20",
        1427 => x"256c750d",
        1428 => x"0a000000",
        1429 => x"232d302b",
        1430 => x"20000000",
        1431 => x"686c4c00",
        1432 => x"65666745",
        1433 => x"46470000",
        1434 => x"30313233",
        1435 => x"34353637",
        1436 => x"38394142",
        1437 => x"43444546",
        1438 => x"00000000",
        1439 => x"30313233",
        1440 => x"34353637",
        1441 => x"38396162",
        1442 => x"63646566",
        1443 => x"00000000",
        1444 => x"180d0000",
        1445 => x"380d0000",
        1446 => x"e40c0000",
        1447 => x"e40c0000",
        1448 => x"e40c0000",
        1449 => x"e40c0000",
        1450 => x"380d0000",
        1451 => x"e40c0000",
        1452 => x"e40c0000",
        1453 => x"e40c0000",
        1454 => x"e40c0000",
        1455 => x"500f0000",
        1456 => x"cc0d0000",
        1457 => x"b80e0000",
        1458 => x"e40c0000",
        1459 => x"e40c0000",
        1460 => x"980f0000",
        1461 => x"e40c0000",
        1462 => x"cc0d0000",
        1463 => x"e40c0000",
        1464 => x"e40c0000",
        1465 => x"c40e0000",
        1466 => x"18000020",
        1467 => x"a4150000",
        1468 => x"ac150000",
        1469 => x"d8150000",
        1470 => x"04160000",
        1471 => x"2c160000",
        1472 => x"00000000",
        1473 => x"00000000",
        1474 => x"00000000",
        1475 => x"00000000",
        1476 => x"00000000",
        1477 => x"00000000",
        1478 => x"00000000",
        1479 => x"00000000",
        1480 => x"00000000",
        1481 => x"00000000",
        1482 => x"00000000",
        1483 => x"00000000",
        1484 => x"00000000",
        1485 => x"00000000",
        1486 => x"00000000",
        1487 => x"00000000",
        1488 => x"00000000",
        1489 => x"00000000",
        1490 => x"00000000",
        1491 => x"00000000",
        1492 => x"00000000",
        1493 => x"00000000",
        1494 => x"00000000",
        1495 => x"00000000",
        1496 => x"00000000",
        1497 => x"18000020",
        others => (others => '0')
    );
end package processor_common_rom;
