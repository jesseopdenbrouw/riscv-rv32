-- srec2vhdl table generator
-- for input file interrupt_direct.srec

library ieee;
use ieee.std_logic_1164.all;

library work;
use work.processor_common.all;

package processor_common_rom is
    constant rom_contents : rom_type := (
           0 => x"97110020",
           1 => x"93810180",
           2 => x"17810020",
           3 => x"130181ff",
           4 => x"97020000",
           5 => x"9382421d",
           6 => x"73905230",
           7 => x"13860188",
           8 => x"93874189",
           9 => x"637af600",
          10 => x"3386c740",
          11 => x"93050000",
          12 => x"13850188",
          13 => x"ef10c049",
          14 => x"37050020",
          15 => x"13060500",
          16 => x"93870188",
          17 => x"637cf600",
          18 => x"b7350000",
          19 => x"3386c740",
          20 => x"93854512",
          21 => x"13050500",
          22 => x"ef104045",
          23 => x"ef105001",
          24 => x"b7050020",
          25 => x"13060000",
          26 => x"93850500",
          27 => x"13055000",
          28 => x"ef10804b",
          29 => x"ef10c07b",
          30 => x"37350000",
          31 => x"130101ff",
          32 => x"130505f7",
          33 => x"23261100",
          34 => x"23248100",
          35 => x"23229100",
          36 => x"23202101",
          37 => x"ef004018",
          38 => x"73294034",
          39 => x"93040002",
          40 => x"37040080",
          41 => x"33758900",
          42 => x"3335a000",
          43 => x"13050503",
          44 => x"9384f4ff",
          45 => x"ef004014",
          46 => x"13541400",
          47 => x"e39404fe",
          48 => x"03248100",
          49 => x"8320c100",
          50 => x"83244100",
          51 => x"03290100",
          52 => x"37350000",
          53 => x"130505fb",
          54 => x"13010101",
          55 => x"6f00c013",
          56 => x"b70700f0",
          57 => x"03a74708",
          58 => x"1377f7fe",
          59 => x"23a2e708",
          60 => x"03a74700",
          61 => x"13471700",
          62 => x"23a2e700",
          63 => x"67800000",
          64 => x"370700f0",
          65 => x"83274700",
          66 => x"93e70720",
          67 => x"2322f700",
          68 => x"6f000000",
          69 => x"b70700f0",
          70 => x"83a6470f",
          71 => x"03a6070f",
          72 => x"03a7470f",
          73 => x"e31ad7fe",
          74 => x"b7860100",
          75 => x"9305f0ff",
          76 => x"9386066a",
          77 => x"23aeb70e",
          78 => x"b306d600",
          79 => x"23acb70e",
          80 => x"33b6c600",
          81 => x"23acd70e",
          82 => x"3306e600",
          83 => x"23aec70e",
          84 => x"03a74700",
          85 => x"13472700",
          86 => x"23a2e700",
          87 => x"67800000",
          88 => x"370700f0",
          89 => x"8327c702",
          90 => x"93f74700",
          91 => x"638a0700",
          92 => x"83274700",
          93 => x"93c78700",
          94 => x"2322f700",
          95 => x"83270702",
          96 => x"67800000",
          97 => x"b70700f0",
          98 => x"03a7470a",
          99 => x"1377f7f0",
         100 => x"23a2e70a",
         101 => x"03a74700",
         102 => x"13474700",
         103 => x"23a2e700",
         104 => x"67800000",
         105 => x"b70700f0",
         106 => x"03a74706",
         107 => x"137777ff",
         108 => x"23a2e706",
         109 => x"03a74700",
         110 => x"13470701",
         111 => x"23a2e700",
         112 => x"67800000",
         113 => x"b70700f0",
         114 => x"03a74704",
         115 => x"137777fe",
         116 => x"23a2e704",
         117 => x"03a74700",
         118 => x"13470702",
         119 => x"23a2e700",
         120 => x"67800000",
         121 => x"6f000000",
         122 => x"b70700f0",
         123 => x"23a2a702",
         124 => x"23a4b702",
         125 => x"67800000",
         126 => x"1375f50f",
         127 => x"b70700f0",
         128 => x"23a0a702",
         129 => x"370700f0",
         130 => x"8327c702",
         131 => x"93f70701",
         132 => x"e38c07fe",
         133 => x"67800000",
         134 => x"63060502",
         135 => x"83470500",
         136 => x"63820702",
         137 => x"370700f0",
         138 => x"13051500",
         139 => x"2320f702",
         140 => x"8327c702",
         141 => x"93f70701",
         142 => x"e38c07fe",
         143 => x"83470500",
         144 => x"e39407fe",
         145 => x"67800000",
         146 => x"370700f0",
         147 => x"8327c702",
         148 => x"93f74700",
         149 => x"e38c07fe",
         150 => x"03250702",
         151 => x"1375f50f",
         152 => x"67800000",
         153 => x"b70700f0",
         154 => x"03a5c702",
         155 => x"13754500",
         156 => x"67800000",
         157 => x"373e0000",
         158 => x"930e0500",
         159 => x"138ff5ff",
         160 => x"13050000",
         161 => x"130e0ed1",
         162 => x"b70600f0",
         163 => x"13035001",
         164 => x"9308f007",
         165 => x"13082000",
         166 => x"93052001",
         167 => x"83a7c602",
         168 => x"93f74700",
         169 => x"e38c07fe",
         170 => x"03a60602",
         171 => x"1377f60f",
         172 => x"6360e302",
         173 => x"6370e802",
         174 => x"9307d7ff",
         175 => x"63ecf500",
         176 => x"93972700",
         177 => x"b307fe00",
         178 => x"83a70700",
         179 => x"67800700",
         180 => x"630e1707",
         181 => x"6352e513",
         182 => x"1376f60f",
         183 => x"930706fe",
         184 => x"93f7f70f",
         185 => x"930fe005",
         186 => x"e3eafffa",
         187 => x"b387ae00",
         188 => x"2380c700",
         189 => x"b70700f0",
         190 => x"23a0e702",
         191 => x"13051500",
         192 => x"370700f0",
         193 => x"8327c702",
         194 => x"93f70701",
         195 => x"e38c07fe",
         196 => x"6ff0dff8",
         197 => x"b38eae00",
         198 => x"b7360000",
         199 => x"23800e00",
         200 => x"9307d000",
         201 => x"938606fb",
         202 => x"370700f0",
         203 => x"93861600",
         204 => x"2320f702",
         205 => x"8327c702",
         206 => x"93f70701",
         207 => x"e38c07fe",
         208 => x"83c70600",
         209 => x"e39407fe",
         210 => x"67800000",
         211 => x"b70700f0",
         212 => x"63040508",
         213 => x"1307f007",
         214 => x"23a0e702",
         215 => x"370700f0",
         216 => x"8327c702",
         217 => x"93f70701",
         218 => x"e38c07fe",
         219 => x"1305f5ff",
         220 => x"6ff0dff2",
         221 => x"370700f0",
         222 => x"13070702",
         223 => x"1306f007",
         224 => x"630e0500",
         225 => x"2320c700",
         226 => x"8327c700",
         227 => x"93f70701",
         228 => x"e38c07fe",
         229 => x"1305f5ff",
         230 => x"e31605fe",
         231 => x"13050000",
         232 => x"6ff0dfef",
         233 => x"37360000",
         234 => x"9307c003",
         235 => x"13060608",
         236 => x"370700f0",
         237 => x"13061600",
         238 => x"2320f702",
         239 => x"8327c702",
         240 => x"93f70701",
         241 => x"e38c07fe",
         242 => x"83470600",
         243 => x"e39407fe",
         244 => x"13050000",
         245 => x"6ff09fec",
         246 => x"13077000",
         247 => x"23a0e702",
         248 => x"370700f0",
         249 => x"8327c702",
         250 => x"93f70701",
         251 => x"e38c07fe",
         252 => x"13050000",
         253 => x"6ff09fea",
         254 => x"13077000",
         255 => x"b70700f0",
         256 => x"23a0e702",
         257 => x"370700f0",
         258 => x"8327c702",
         259 => x"93f70701",
         260 => x"e38c07fe",
         261 => x"6ff09fe8",
         262 => x"1375f50f",
         263 => x"b70700f0",
         264 => x"23a0a702",
         265 => x"370700f0",
         266 => x"8327c702",
         267 => x"93f70701",
         268 => x"e38c07fe",
         269 => x"13051000",
         270 => x"67800000",
         271 => x"370700f0",
         272 => x"8327c702",
         273 => x"93f74700",
         274 => x"e38c07fe",
         275 => x"03250702",
         276 => x"1375f50f",
         277 => x"67800000",
         278 => x"13050000",
         279 => x"67800000",
         280 => x"13050000",
         281 => x"67800000",
         282 => x"130101f8",
         283 => x"23221100",
         284 => x"23242100",
         285 => x"23263100",
         286 => x"23284100",
         287 => x"232a5100",
         288 => x"232c6100",
         289 => x"232e7100",
         290 => x"23208102",
         291 => x"23229102",
         292 => x"2324a102",
         293 => x"2326b102",
         294 => x"2328c102",
         295 => x"232ad102",
         296 => x"232ce102",
         297 => x"232ef102",
         298 => x"23200105",
         299 => x"23221105",
         300 => x"23242105",
         301 => x"23263105",
         302 => x"23284105",
         303 => x"232a5105",
         304 => x"232c6105",
         305 => x"232e7105",
         306 => x"23208107",
         307 => x"23229107",
         308 => x"2324a107",
         309 => x"2326b107",
         310 => x"2328c107",
         311 => x"232ad107",
         312 => x"232ce107",
         313 => x"232ef107",
         314 => x"f3272034",
         315 => x"37070080",
         316 => x"93067700",
         317 => x"6386d70e",
         318 => x"9306b000",
         319 => x"63fef602",
         320 => x"9346f7fe",
         321 => x"b386d700",
         322 => x"13064000",
         323 => x"636ad602",
         324 => x"1347e7fe",
         325 => x"b387e700",
         326 => x"13073000",
         327 => x"6364f714",
         328 => x"37370000",
         329 => x"93972700",
         330 => x"1307c7d5",
         331 => x"b387e700",
         332 => x"83a70700",
         333 => x"67800700",
         334 => x"13071000",
         335 => x"6364f708",
         336 => x"03258102",
         337 => x"832fc107",
         338 => x"032f8107",
         339 => x"832e4107",
         340 => x"032e0107",
         341 => x"832dc106",
         342 => x"032d8106",
         343 => x"832c4106",
         344 => x"032c0106",
         345 => x"832bc105",
         346 => x"032b8105",
         347 => x"832a4105",
         348 => x"032a0105",
         349 => x"8329c104",
         350 => x"03298104",
         351 => x"83284104",
         352 => x"03280104",
         353 => x"8327c103",
         354 => x"03278103",
         355 => x"83264103",
         356 => x"03260103",
         357 => x"8325c102",
         358 => x"83244102",
         359 => x"03240102",
         360 => x"8323c101",
         361 => x"03238101",
         362 => x"83224101",
         363 => x"03220101",
         364 => x"8321c100",
         365 => x"03218100",
         366 => x"83204100",
         367 => x"13010108",
         368 => x"73002030",
         369 => x"e3eef6f6",
         370 => x"37370000",
         371 => x"93972700",
         372 => x"1307c7d6",
         373 => x"b387e700",
         374 => x"83a70700",
         375 => x"67800700",
         376 => x"eff05fb3",
         377 => x"03258102",
         378 => x"6ff0dff5",
         379 => x"eff09fb9",
         380 => x"03258102",
         381 => x"6ff01ff5",
         382 => x"eff0dfba",
         383 => x"03258102",
         384 => x"6ff05ff4",
         385 => x"eff01fbc",
         386 => x"03258102",
         387 => x"6ff09ff3",
         388 => x"eff01fb5",
         389 => x"03258102",
         390 => x"6ff0dff2",
         391 => x"9307600d",
         392 => x"6384f806",
         393 => x"9307900a",
         394 => x"6388f818",
         395 => x"63ca170f",
         396 => x"938878fc",
         397 => x"93074002",
         398 => x"63ec1703",
         399 => x"b7370000",
         400 => x"9387c7d9",
         401 => x"93982800",
         402 => x"b388f800",
         403 => x"83a70800",
         404 => x"67800700",
         405 => x"13050100",
         406 => x"eff01fa2",
         407 => x"03258102",
         408 => x"6ff05fee",
         409 => x"eff0dfa7",
         410 => x"03258102",
         411 => x"6ff09fed",
         412 => x"ef10801b",
         413 => x"93078005",
         414 => x"2320f500",
         415 => x"9307f0ff",
         416 => x"13850700",
         417 => x"6ff01fec",
         418 => x"63120510",
         419 => x"13858189",
         420 => x"13050500",
         421 => x"6ff01feb",
         422 => x"b7270000",
         423 => x"23a2f500",
         424 => x"93070000",
         425 => x"13850700",
         426 => x"6ff0dfe9",
         427 => x"93070000",
         428 => x"13850700",
         429 => x"6ff01fe9",
         430 => x"ef100017",
         431 => x"93079000",
         432 => x"2320f500",
         433 => x"9307f0ff",
         434 => x"13850700",
         435 => x"6ff09fe7",
         436 => x"13090600",
         437 => x"13840500",
         438 => x"635cc000",
         439 => x"b384c500",
         440 => x"03450400",
         441 => x"13041400",
         442 => x"eff01fd3",
         443 => x"e39a84fe",
         444 => x"13050900",
         445 => x"6ff01fe5",
         446 => x"13090600",
         447 => x"13840500",
         448 => x"e358c0fe",
         449 => x"b384c500",
         450 => x"eff05fd3",
         451 => x"2300a400",
         452 => x"13041400",
         453 => x"e31a94fe",
         454 => x"13050900",
         455 => x"6ff09fe2",
         456 => x"938808c0",
         457 => x"9307f000",
         458 => x"e3e417f5",
         459 => x"b7370000",
         460 => x"938707e3",
         461 => x"93982800",
         462 => x"b388f800",
         463 => x"83a70800",
         464 => x"67800700",
         465 => x"ef10400e",
         466 => x"9307d000",
         467 => x"2320f500",
         468 => x"9307f0ff",
         469 => x"13850700",
         470 => x"6ff0dfde",
         471 => x"ef10c00c",
         472 => x"93072000",
         473 => x"2320f500",
         474 => x"9307f0ff",
         475 => x"13850700",
         476 => x"6ff05fdd",
         477 => x"ef10400b",
         478 => x"9307f001",
         479 => x"2320f500",
         480 => x"9307f0ff",
         481 => x"13850700",
         482 => x"6ff0dfdb",
         483 => x"b7870020",
         484 => x"93870700",
         485 => x"13070040",
         486 => x"b387e740",
         487 => x"e36af5ee",
         488 => x"ef108008",
         489 => x"9307c000",
         490 => x"2320f500",
         491 => x"1305f0ff",
         492 => x"13050500",
         493 => x"6ff01fd9",
         494 => x"13090000",
         495 => x"93040500",
         496 => x"13040900",
         497 => x"93090900",
         498 => x"93070900",
         499 => x"732410c8",
         500 => x"f32910c0",
         501 => x"f32710c8",
         502 => x"e31af4fe",
         503 => x"37460f00",
         504 => x"13060624",
         505 => x"93060000",
         506 => x"13850900",
         507 => x"93050400",
         508 => x"ef00900d",
         509 => x"37460f00",
         510 => x"23a4a400",
         511 => x"13060624",
         512 => x"93060000",
         513 => x"13850900",
         514 => x"93050400",
         515 => x"ef00c048",
         516 => x"23a0a400",
         517 => x"23a2b400",
         518 => x"13050900",
         519 => x"6ff09fd2",
         520 => x"13030500",
         521 => x"138e0500",
         522 => x"93080000",
         523 => x"63dc0500",
         524 => x"b337a000",
         525 => x"330eb040",
         526 => x"330efe40",
         527 => x"3303a040",
         528 => x"9308f0ff",
         529 => x"63dc0600",
         530 => x"b337c000",
         531 => x"b306d040",
         532 => x"93c8f8ff",
         533 => x"b386f640",
         534 => x"3306c040",
         535 => x"13070600",
         536 => x"13080300",
         537 => x"93070e00",
         538 => x"639c0628",
         539 => x"b7350000",
         540 => x"938505e7",
         541 => x"6376ce0e",
         542 => x"b7060100",
         543 => x"6378d60c",
         544 => x"93360610",
         545 => x"93c61600",
         546 => x"93963600",
         547 => x"3355d600",
         548 => x"b385a500",
         549 => x"83c50500",
         550 => x"13050002",
         551 => x"b386d500",
         552 => x"b305d540",
         553 => x"630cd500",
         554 => x"b317be00",
         555 => x"b356d300",
         556 => x"3317b600",
         557 => x"b3e7f600",
         558 => x"3318b300",
         559 => x"93550701",
         560 => x"33deb702",
         561 => x"13160701",
         562 => x"13560601",
         563 => x"b3f7b702",
         564 => x"13050e00",
         565 => x"3303c603",
         566 => x"93960701",
         567 => x"93570801",
         568 => x"b3e7d700",
         569 => x"63fe6700",
         570 => x"b307f700",
         571 => x"1305feff",
         572 => x"63e8e700",
         573 => x"63f66700",
         574 => x"1305eeff",
         575 => x"b387e700",
         576 => x"b3876740",
         577 => x"33d3b702",
         578 => x"13180801",
         579 => x"13580801",
         580 => x"b3f7b702",
         581 => x"b3066602",
         582 => x"93970701",
         583 => x"3368f800",
         584 => x"93070300",
         585 => x"637cd800",
         586 => x"33080701",
         587 => x"9307f3ff",
         588 => x"6366e800",
         589 => x"6374d800",
         590 => x"9307e3ff",
         591 => x"13150501",
         592 => x"3365f500",
         593 => x"93050000",
         594 => x"6f00000e",
         595 => x"37050001",
         596 => x"93060001",
         597 => x"e36ca6f2",
         598 => x"93068001",
         599 => x"6ff01ff3",
         600 => x"93060000",
         601 => x"630c0600",
         602 => x"b7070100",
         603 => x"637af60c",
         604 => x"93360610",
         605 => x"93c61600",
         606 => x"93963600",
         607 => x"b357d600",
         608 => x"b385f500",
         609 => x"83c70500",
         610 => x"b387d700",
         611 => x"93060002",
         612 => x"b385f640",
         613 => x"6390f60c",
         614 => x"b307ce40",
         615 => x"93051000",
         616 => x"13530701",
         617 => x"b3de6702",
         618 => x"13160701",
         619 => x"13560601",
         620 => x"93560801",
         621 => x"b3f76702",
         622 => x"13850e00",
         623 => x"330ed603",
         624 => x"93970701",
         625 => x"b3e7f600",
         626 => x"63fec701",
         627 => x"b307f700",
         628 => x"1385feff",
         629 => x"63e8e700",
         630 => x"63f6c701",
         631 => x"1385eeff",
         632 => x"b387e700",
         633 => x"b387c741",
         634 => x"33de6702",
         635 => x"13180801",
         636 => x"13580801",
         637 => x"b3f76702",
         638 => x"b306c603",
         639 => x"93970701",
         640 => x"3368f800",
         641 => x"93070e00",
         642 => x"637cd800",
         643 => x"33080701",
         644 => x"9307feff",
         645 => x"6366e800",
         646 => x"6374d800",
         647 => x"9307eeff",
         648 => x"13150501",
         649 => x"3365f500",
         650 => x"638a0800",
         651 => x"b337a000",
         652 => x"b305b040",
         653 => x"b385f540",
         654 => x"3305a040",
         655 => x"67800000",
         656 => x"b7070001",
         657 => x"93060001",
         658 => x"e36af6f2",
         659 => x"93068001",
         660 => x"6ff0dff2",
         661 => x"3317b600",
         662 => x"b356fe00",
         663 => x"13550701",
         664 => x"331ebe00",
         665 => x"b357f300",
         666 => x"b3e7c701",
         667 => x"33dea602",
         668 => x"13160701",
         669 => x"13560601",
         670 => x"3318b300",
         671 => x"b3f6a602",
         672 => x"3303c603",
         673 => x"93950601",
         674 => x"93d60701",
         675 => x"b3e6b600",
         676 => x"93050e00",
         677 => x"63fe6600",
         678 => x"b306d700",
         679 => x"9305feff",
         680 => x"63e8e600",
         681 => x"63f66600",
         682 => x"9305eeff",
         683 => x"b386e600",
         684 => x"b3866640",
         685 => x"33d3a602",
         686 => x"93970701",
         687 => x"93d70701",
         688 => x"b3f6a602",
         689 => x"33066602",
         690 => x"93960601",
         691 => x"b3e7d700",
         692 => x"93060300",
         693 => x"63fec700",
         694 => x"b307f700",
         695 => x"9306f3ff",
         696 => x"63e8e700",
         697 => x"63f6c700",
         698 => x"9306e3ff",
         699 => x"b387e700",
         700 => x"93950501",
         701 => x"b387c740",
         702 => x"b3e5d500",
         703 => x"6ff05fea",
         704 => x"6366de18",
         705 => x"b7070100",
         706 => x"63f4f604",
         707 => x"13b70610",
         708 => x"13471700",
         709 => x"13173700",
         710 => x"b7370000",
         711 => x"b3d5e600",
         712 => x"938707e7",
         713 => x"b387b700",
         714 => x"83c70700",
         715 => x"b387e700",
         716 => x"13070002",
         717 => x"b305f740",
         718 => x"6316f702",
         719 => x"13051000",
         720 => x"e3e4c6ef",
         721 => x"3335c300",
         722 => x"13451500",
         723 => x"6ff0dfed",
         724 => x"b7070001",
         725 => x"13070001",
         726 => x"e3e0f6fc",
         727 => x"13078001",
         728 => x"6ff09ffb",
         729 => x"3357f600",
         730 => x"b396b600",
         731 => x"b366d700",
         732 => x"3357fe00",
         733 => x"331ebe00",
         734 => x"b357f300",
         735 => x"b3e7c701",
         736 => x"13de0601",
         737 => x"335fc703",
         738 => x"13980601",
         739 => x"13580801",
         740 => x"3316b600",
         741 => x"3377c703",
         742 => x"b30ee803",
         743 => x"13150701",
         744 => x"13d70701",
         745 => x"3367a700",
         746 => x"13050f00",
         747 => x"637ed701",
         748 => x"3387e600",
         749 => x"1305ffff",
         750 => x"6368d700",
         751 => x"6376d701",
         752 => x"1305efff",
         753 => x"3307d700",
         754 => x"3307d741",
         755 => x"b35ec703",
         756 => x"93970701",
         757 => x"93d70701",
         758 => x"3377c703",
         759 => x"3308d803",
         760 => x"13170701",
         761 => x"b3e7e700",
         762 => x"13870e00",
         763 => x"63fe0701",
         764 => x"b387f600",
         765 => x"1387feff",
         766 => x"63e8d700",
         767 => x"63f60701",
         768 => x"1387eeff",
         769 => x"b387d700",
         770 => x"13150501",
         771 => x"b70e0100",
         772 => x"3365e500",
         773 => x"9386feff",
         774 => x"3377d500",
         775 => x"b3870741",
         776 => x"b376d600",
         777 => x"13580501",
         778 => x"13560601",
         779 => x"330ed702",
         780 => x"b306d802",
         781 => x"3307c702",
         782 => x"3308c802",
         783 => x"3306d700",
         784 => x"13570e01",
         785 => x"3307c700",
         786 => x"6374d700",
         787 => x"3308d801",
         788 => x"93560701",
         789 => x"b3860601",
         790 => x"63e6d702",
         791 => x"e394d7ce",
         792 => x"b7070100",
         793 => x"9387f7ff",
         794 => x"3377f700",
         795 => x"13170701",
         796 => x"337efe00",
         797 => x"3313b300",
         798 => x"3307c701",
         799 => x"93050000",
         800 => x"e374e3da",
         801 => x"1305f5ff",
         802 => x"6ff0dfcb",
         803 => x"93050000",
         804 => x"13050000",
         805 => x"6ff05fd9",
         806 => x"93080500",
         807 => x"13830500",
         808 => x"13070600",
         809 => x"13080500",
         810 => x"93870500",
         811 => x"63920628",
         812 => x"b7350000",
         813 => x"938505e7",
         814 => x"6376c30e",
         815 => x"b7060100",
         816 => x"6378d60c",
         817 => x"93360610",
         818 => x"93c61600",
         819 => x"93963600",
         820 => x"3355d600",
         821 => x"b385a500",
         822 => x"83c50500",
         823 => x"13050002",
         824 => x"b386d500",
         825 => x"b305d540",
         826 => x"630cd500",
         827 => x"b317b300",
         828 => x"b3d6d800",
         829 => x"3317b600",
         830 => x"b3e7f600",
         831 => x"3398b800",
         832 => x"93550701",
         833 => x"33d3b702",
         834 => x"13160701",
         835 => x"13560601",
         836 => x"b3f7b702",
         837 => x"13050300",
         838 => x"b3086602",
         839 => x"93960701",
         840 => x"93570801",
         841 => x"b3e7d700",
         842 => x"63fe1701",
         843 => x"b307f700",
         844 => x"1305f3ff",
         845 => x"63e8e700",
         846 => x"63f61701",
         847 => x"1305e3ff",
         848 => x"b387e700",
         849 => x"b3871741",
         850 => x"b3d8b702",
         851 => x"13180801",
         852 => x"13580801",
         853 => x"b3f7b702",
         854 => x"b3061603",
         855 => x"93970701",
         856 => x"3368f800",
         857 => x"93870800",
         858 => x"637cd800",
         859 => x"33080701",
         860 => x"9387f8ff",
         861 => x"6366e800",
         862 => x"6374d800",
         863 => x"9387e8ff",
         864 => x"13150501",
         865 => x"3365f500",
         866 => x"93050000",
         867 => x"67800000",
         868 => x"37050001",
         869 => x"93060001",
         870 => x"e36ca6f2",
         871 => x"93068001",
         872 => x"6ff01ff3",
         873 => x"93060000",
         874 => x"630c0600",
         875 => x"b7070100",
         876 => x"6370f60c",
         877 => x"93360610",
         878 => x"93c61600",
         879 => x"93963600",
         880 => x"b357d600",
         881 => x"b385f500",
         882 => x"83c70500",
         883 => x"b387d700",
         884 => x"93060002",
         885 => x"b385f640",
         886 => x"6396f60a",
         887 => x"b307c340",
         888 => x"93051000",
         889 => x"93580701",
         890 => x"33de1703",
         891 => x"13160701",
         892 => x"13560601",
         893 => x"93560801",
         894 => x"b3f71703",
         895 => x"13050e00",
         896 => x"3303c603",
         897 => x"93970701",
         898 => x"b3e7f600",
         899 => x"63fe6700",
         900 => x"b307f700",
         901 => x"1305feff",
         902 => x"63e8e700",
         903 => x"63f66700",
         904 => x"1305eeff",
         905 => x"b387e700",
         906 => x"b3876740",
         907 => x"33d31703",
         908 => x"13180801",
         909 => x"13580801",
         910 => x"b3f71703",
         911 => x"b3066602",
         912 => x"93970701",
         913 => x"3368f800",
         914 => x"93070300",
         915 => x"637cd800",
         916 => x"33080701",
         917 => x"9307f3ff",
         918 => x"6366e800",
         919 => x"6374d800",
         920 => x"9307e3ff",
         921 => x"13150501",
         922 => x"3365f500",
         923 => x"67800000",
         924 => x"b7070001",
         925 => x"93060001",
         926 => x"e364f6f4",
         927 => x"93068001",
         928 => x"6ff01ff4",
         929 => x"3317b600",
         930 => x"b356f300",
         931 => x"13550701",
         932 => x"3313b300",
         933 => x"b3d7f800",
         934 => x"b3e76700",
         935 => x"33d3a602",
         936 => x"13160701",
         937 => x"13560601",
         938 => x"3398b800",
         939 => x"b3f6a602",
         940 => x"b3086602",
         941 => x"93950601",
         942 => x"93d60701",
         943 => x"b3e6b600",
         944 => x"93050300",
         945 => x"63fe1601",
         946 => x"b306d700",
         947 => x"9305f3ff",
         948 => x"63e8e600",
         949 => x"63f61601",
         950 => x"9305e3ff",
         951 => x"b386e600",
         952 => x"b3861641",
         953 => x"b3d8a602",
         954 => x"93970701",
         955 => x"93d70701",
         956 => x"b3f6a602",
         957 => x"33061603",
         958 => x"93960601",
         959 => x"b3e7d700",
         960 => x"93860800",
         961 => x"63fec700",
         962 => x"b307f700",
         963 => x"9386f8ff",
         964 => x"63e8e700",
         965 => x"63f6c700",
         966 => x"9386e8ff",
         967 => x"b387e700",
         968 => x"93950501",
         969 => x"b387c740",
         970 => x"b3e5d500",
         971 => x"6ff09feb",
         972 => x"63e6d518",
         973 => x"b7070100",
         974 => x"63f4f604",
         975 => x"13b70610",
         976 => x"13471700",
         977 => x"13173700",
         978 => x"b7370000",
         979 => x"b3d5e600",
         980 => x"938707e7",
         981 => x"b387b700",
         982 => x"83c70700",
         983 => x"b387e700",
         984 => x"13070002",
         985 => x"b305f740",
         986 => x"6316f702",
         987 => x"13051000",
         988 => x"e3ee66e0",
         989 => x"33b5c800",
         990 => x"13451500",
         991 => x"67800000",
         992 => x"b7070001",
         993 => x"13070001",
         994 => x"e3e0f6fc",
         995 => x"13078001",
         996 => x"6ff09ffb",
         997 => x"3357f600",
         998 => x"b396b600",
         999 => x"b366d700",
        1000 => x"3357f300",
        1001 => x"3313b300",
        1002 => x"b3d7f800",
        1003 => x"b3e76700",
        1004 => x"13d30601",
        1005 => x"b35e6702",
        1006 => x"13980601",
        1007 => x"13580801",
        1008 => x"3316b600",
        1009 => x"33776702",
        1010 => x"330ed803",
        1011 => x"13150701",
        1012 => x"13d70701",
        1013 => x"3367a700",
        1014 => x"13850e00",
        1015 => x"637ec701",
        1016 => x"3387e600",
        1017 => x"1385feff",
        1018 => x"6368d700",
        1019 => x"6376c701",
        1020 => x"1385eeff",
        1021 => x"3307d700",
        1022 => x"3307c741",
        1023 => x"335e6702",
        1024 => x"93970701",
        1025 => x"93d70701",
        1026 => x"33776702",
        1027 => x"3308c803",
        1028 => x"13170701",
        1029 => x"b3e7e700",
        1030 => x"13070e00",
        1031 => x"63fe0701",
        1032 => x"b387f600",
        1033 => x"1307feff",
        1034 => x"63e8d700",
        1035 => x"63f60701",
        1036 => x"1307eeff",
        1037 => x"b387d700",
        1038 => x"13150501",
        1039 => x"370e0100",
        1040 => x"3365e500",
        1041 => x"9306feff",
        1042 => x"3377d500",
        1043 => x"b3870741",
        1044 => x"b376d600",
        1045 => x"13580501",
        1046 => x"13560601",
        1047 => x"3303d702",
        1048 => x"b306d802",
        1049 => x"3307c702",
        1050 => x"3308c802",
        1051 => x"3306d700",
        1052 => x"13570301",
        1053 => x"3307c700",
        1054 => x"6374d700",
        1055 => x"3308c801",
        1056 => x"93560701",
        1057 => x"b3860601",
        1058 => x"63e6d702",
        1059 => x"e39ed7ce",
        1060 => x"b7070100",
        1061 => x"9387f7ff",
        1062 => x"3377f700",
        1063 => x"13170701",
        1064 => x"3373f300",
        1065 => x"b398b800",
        1066 => x"33076700",
        1067 => x"93050000",
        1068 => x"e3fee8cc",
        1069 => x"1305f5ff",
        1070 => x"6ff01fcd",
        1071 => x"93050000",
        1072 => x"13050000",
        1073 => x"67800000",
        1074 => x"13080600",
        1075 => x"93070500",
        1076 => x"13870500",
        1077 => x"63960620",
        1078 => x"b7380000",
        1079 => x"938808e7",
        1080 => x"63fcc50c",
        1081 => x"b7060100",
        1082 => x"637ed60a",
        1083 => x"93360610",
        1084 => x"93c61600",
        1085 => x"93963600",
        1086 => x"3353d600",
        1087 => x"b3886800",
        1088 => x"83c80800",
        1089 => x"13030002",
        1090 => x"b386d800",
        1091 => x"b308d340",
        1092 => x"630cd300",
        1093 => x"33971501",
        1094 => x"b356d500",
        1095 => x"33181601",
        1096 => x"33e7e600",
        1097 => x"b3171501",
        1098 => x"13560801",
        1099 => x"b356c702",
        1100 => x"13150801",
        1101 => x"13550501",
        1102 => x"3377c702",
        1103 => x"b386a602",
        1104 => x"93150701",
        1105 => x"13d70701",
        1106 => x"3367b700",
        1107 => x"637ad700",
        1108 => x"3307e800",
        1109 => x"63660701",
        1110 => x"6374d700",
        1111 => x"33070701",
        1112 => x"3307d740",
        1113 => x"b356c702",
        1114 => x"3377c702",
        1115 => x"b386a602",
        1116 => x"93970701",
        1117 => x"13170701",
        1118 => x"93d70701",
        1119 => x"b3e7e700",
        1120 => x"63fad700",
        1121 => x"b307f800",
        1122 => x"63e60701",
        1123 => x"63f4d700",
        1124 => x"b3870701",
        1125 => x"b387d740",
        1126 => x"33d51701",
        1127 => x"93050000",
        1128 => x"67800000",
        1129 => x"37030001",
        1130 => x"93060001",
        1131 => x"e36666f4",
        1132 => x"93068001",
        1133 => x"6ff05ff4",
        1134 => x"93060000",
        1135 => x"630c0600",
        1136 => x"37070100",
        1137 => x"637ee606",
        1138 => x"93360610",
        1139 => x"93c61600",
        1140 => x"93963600",
        1141 => x"3357d600",
        1142 => x"b388e800",
        1143 => x"03c70800",
        1144 => x"3307d700",
        1145 => x"93060002",
        1146 => x"b388e640",
        1147 => x"6394e606",
        1148 => x"3387c540",
        1149 => x"93550801",
        1150 => x"3356b702",
        1151 => x"13150801",
        1152 => x"13550501",
        1153 => x"93d60701",
        1154 => x"3377b702",
        1155 => x"3306a602",
        1156 => x"13170701",
        1157 => x"33e7e600",
        1158 => x"637ac700",
        1159 => x"3307e800",
        1160 => x"63660701",
        1161 => x"6374c700",
        1162 => x"33070701",
        1163 => x"3307c740",
        1164 => x"b356b702",
        1165 => x"3377b702",
        1166 => x"b386a602",
        1167 => x"6ff05ff3",
        1168 => x"37070001",
        1169 => x"93060001",
        1170 => x"e366e6f8",
        1171 => x"93068001",
        1172 => x"6ff05ff8",
        1173 => x"33181601",
        1174 => x"b3d6e500",
        1175 => x"b3171501",
        1176 => x"b3951501",
        1177 => x"3357e500",
        1178 => x"13550801",
        1179 => x"3367b700",
        1180 => x"b3d5a602",
        1181 => x"13130801",
        1182 => x"13530301",
        1183 => x"b3f6a602",
        1184 => x"b3856502",
        1185 => x"13960601",
        1186 => x"93560701",
        1187 => x"b3e6c600",
        1188 => x"63fab600",
        1189 => x"b306d800",
        1190 => x"63e60601",
        1191 => x"63f4b600",
        1192 => x"b3860601",
        1193 => x"b386b640",
        1194 => x"33d6a602",
        1195 => x"13170701",
        1196 => x"13570701",
        1197 => x"b3f6a602",
        1198 => x"33066602",
        1199 => x"93960601",
        1200 => x"3367d700",
        1201 => x"637ac700",
        1202 => x"3307e800",
        1203 => x"63660701",
        1204 => x"6374c700",
        1205 => x"33070701",
        1206 => x"3307c740",
        1207 => x"6ff09ff1",
        1208 => x"63e4d51c",
        1209 => x"37080100",
        1210 => x"63fe0605",
        1211 => x"13b80610",
        1212 => x"13481800",
        1213 => x"13183800",
        1214 => x"b7380000",
        1215 => x"33d30601",
        1216 => x"938808e7",
        1217 => x"b3886800",
        1218 => x"83c80800",
        1219 => x"13030002",
        1220 => x"b3880801",
        1221 => x"33081341",
        1222 => x"63101305",
        1223 => x"63e4b600",
        1224 => x"636cc500",
        1225 => x"3306c540",
        1226 => x"b386d540",
        1227 => x"3337c500",
        1228 => x"93070600",
        1229 => x"3387e640",
        1230 => x"13850700",
        1231 => x"93050700",
        1232 => x"67800000",
        1233 => x"b7080001",
        1234 => x"13080001",
        1235 => x"e3e616fb",
        1236 => x"13088001",
        1237 => x"6ff05ffa",
        1238 => x"b3571601",
        1239 => x"b3960601",
        1240 => x"b3e6d700",
        1241 => x"33d71501",
        1242 => x"13de0601",
        1243 => x"335fc703",
        1244 => x"13930601",
        1245 => x"13530301",
        1246 => x"b3970501",
        1247 => x"b3551501",
        1248 => x"b3e5f500",
        1249 => x"93d70501",
        1250 => x"33160601",
        1251 => x"33150501",
        1252 => x"3377c703",
        1253 => x"b30ee303",
        1254 => x"13170701",
        1255 => x"b3e7e700",
        1256 => x"13070f00",
        1257 => x"63fed701",
        1258 => x"b387f600",
        1259 => x"1307ffff",
        1260 => x"63e8d700",
        1261 => x"63f6d701",
        1262 => x"1307efff",
        1263 => x"b387d700",
        1264 => x"b387d741",
        1265 => x"b3dec703",
        1266 => x"93950501",
        1267 => x"93d50501",
        1268 => x"b3f7c703",
        1269 => x"138e0e00",
        1270 => x"3303d303",
        1271 => x"93970701",
        1272 => x"b3e5f500",
        1273 => x"63fe6500",
        1274 => x"b385b600",
        1275 => x"138efeff",
        1276 => x"63e8d500",
        1277 => x"63f66500",
        1278 => x"138eeeff",
        1279 => x"b385d500",
        1280 => x"93170701",
        1281 => x"370f0100",
        1282 => x"b3e7c701",
        1283 => x"b3856540",
        1284 => x"1303ffff",
        1285 => x"33f76700",
        1286 => x"135e0601",
        1287 => x"93d70701",
        1288 => x"33736600",
        1289 => x"b30e6702",
        1290 => x"33836702",
        1291 => x"3307c703",
        1292 => x"b387c703",
        1293 => x"330e6700",
        1294 => x"13d70e01",
        1295 => x"3307c701",
        1296 => x"63746700",
        1297 => x"b387e701",
        1298 => x"13530701",
        1299 => x"b307f300",
        1300 => x"37030100",
        1301 => x"1303f3ff",
        1302 => x"33776700",
        1303 => x"13170701",
        1304 => x"b3fe6e00",
        1305 => x"3307d701",
        1306 => x"63e6f500",
        1307 => x"639ef500",
        1308 => x"637ce500",
        1309 => x"3306c740",
        1310 => x"3333c700",
        1311 => x"b306d300",
        1312 => x"13070600",
        1313 => x"b387d740",
        1314 => x"3307e540",
        1315 => x"3335e500",
        1316 => x"b385f540",
        1317 => x"b385a540",
        1318 => x"b3981501",
        1319 => x"33570701",
        1320 => x"33e5e800",
        1321 => x"b3d50501",
        1322 => x"67800000",
        1323 => x"13030500",
        1324 => x"630e0600",
        1325 => x"83830500",
        1326 => x"23007300",
        1327 => x"1306f6ff",
        1328 => x"13031300",
        1329 => x"93851500",
        1330 => x"e31606fe",
        1331 => x"67800000",
        1332 => x"13030500",
        1333 => x"630a0600",
        1334 => x"2300b300",
        1335 => x"1306f6ff",
        1336 => x"13031300",
        1337 => x"e31a06fe",
        1338 => x"67800000",
        1339 => x"630c0602",
        1340 => x"13030500",
        1341 => x"93061000",
        1342 => x"636ab500",
        1343 => x"9306f0ff",
        1344 => x"1307f6ff",
        1345 => x"3303e300",
        1346 => x"b385e500",
        1347 => x"83830500",
        1348 => x"23007300",
        1349 => x"1306f6ff",
        1350 => x"3303d300",
        1351 => x"b385d500",
        1352 => x"e31606fe",
        1353 => x"67800000",
        1354 => x"130101f9",
        1355 => x"23248106",
        1356 => x"23229106",
        1357 => x"23261106",
        1358 => x"23202107",
        1359 => x"232e3105",
        1360 => x"232c4105",
        1361 => x"232a5105",
        1362 => x"23286105",
        1363 => x"23267105",
        1364 => x"23248105",
        1365 => x"23229105",
        1366 => x"2320a105",
        1367 => x"93040500",
        1368 => x"13840500",
        1369 => x"232c0100",
        1370 => x"232e0100",
        1371 => x"23200102",
        1372 => x"23220102",
        1373 => x"23240102",
        1374 => x"23260102",
        1375 => x"23280102",
        1376 => x"232a0102",
        1377 => x"232c0102",
        1378 => x"232e0102",
        1379 => x"97f2ffff",
        1380 => x"9382c2ed",
        1381 => x"73905230",
        1382 => x"93050004",
        1383 => x"1305101b",
        1384 => x"efe09fc4",
        1385 => x"37877d01",
        1386 => x"b70700f0",
        1387 => x"1307f783",
        1388 => x"23a6e708",
        1389 => x"93061001",
        1390 => x"37170000",
        1391 => x"23a0d708",
        1392 => x"13077738",
        1393 => x"23a8e70a",
        1394 => x"37270000",
        1395 => x"1307f770",
        1396 => x"23a6e70a",
        1397 => x"23a0d70a",
        1398 => x"13078070",
        1399 => x"23a0e706",
        1400 => x"3707f900",
        1401 => x"13078700",
        1402 => x"23a0e704",
        1403 => x"93020008",
        1404 => x"73904230",
        1405 => x"b7220000",
        1406 => x"93828280",
        1407 => x"73900230",
        1408 => x"b7390000",
        1409 => x"138509fb",
        1410 => x"efe01fc1",
        1411 => x"63549002",
        1412 => x"1389f4ff",
        1413 => x"9304f0ff",
        1414 => x"03250400",
        1415 => x"1309f9ff",
        1416 => x"13044400",
        1417 => x"efe05fbf",
        1418 => x"138509fb",
        1419 => x"efe0dfbe",
        1420 => x"e31499fe",
        1421 => x"37350000",
        1422 => x"b7faeeee",
        1423 => x"130545f8",
        1424 => x"b7090010",
        1425 => x"37140000",
        1426 => x"1389faee",
        1427 => x"efe0dfbc",
        1428 => x"373b0000",
        1429 => x"9389f9ff",
        1430 => x"938aeaee",
        1431 => x"130404e1",
        1432 => x"93040000",
        1433 => x"b71b0000",
        1434 => x"938b0b2c",
        1435 => x"130af000",
        1436 => x"93050000",
        1437 => x"13058100",
        1438 => x"ef008036",
        1439 => x"938bfbff",
        1440 => x"630a0502",
        1441 => x"e3960bfe",
        1442 => x"73001000",
        1443 => x"b70700f0",
        1444 => x"9306f00f",
        1445 => x"23a4d706",
        1446 => x"03a70704",
        1447 => x"93860704",
        1448 => x"13670730",
        1449 => x"23a0e704",
        1450 => x"93070009",
        1451 => x"23a4f600",
        1452 => x"6ff05ffb",
        1453 => x"032c8100",
        1454 => x"8325c100",
        1455 => x"13060400",
        1456 => x"9357cc01",
        1457 => x"13974500",
        1458 => x"b367f700",
        1459 => x"b3f73701",
        1460 => x"33773c01",
        1461 => x"13d5f541",
        1462 => x"13d88501",
        1463 => x"3307f700",
        1464 => x"33070701",
        1465 => x"9377d500",
        1466 => x"3307f700",
        1467 => x"33774703",
        1468 => x"937725ff",
        1469 => x"93860400",
        1470 => x"13050c00",
        1471 => x"3307f700",
        1472 => x"b307ec40",
        1473 => x"1357f741",
        1474 => x"3338fc00",
        1475 => x"3387e540",
        1476 => x"33070741",
        1477 => x"b3885703",
        1478 => x"33072703",
        1479 => x"33b82703",
        1480 => x"33071701",
        1481 => x"b3872703",
        1482 => x"33070701",
        1483 => x"1358f741",
        1484 => x"13783800",
        1485 => x"b307f800",
        1486 => x"33b80701",
        1487 => x"3307e800",
        1488 => x"1318e701",
        1489 => x"93d72700",
        1490 => x"b367f800",
        1491 => x"13582740",
        1492 => x"93184800",
        1493 => x"13d3c701",
        1494 => x"33e36800",
        1495 => x"33733301",
        1496 => x"b3f83701",
        1497 => x"135e8801",
        1498 => x"1357f741",
        1499 => x"b3886800",
        1500 => x"b388c801",
        1501 => x"1373d700",
        1502 => x"b3886800",
        1503 => x"b3f84803",
        1504 => x"137727ff",
        1505 => x"939c4700",
        1506 => x"b38cfc40",
        1507 => x"939c2c00",
        1508 => x"b30c9c41",
        1509 => x"b388e800",
        1510 => x"33871741",
        1511 => x"93d8f841",
        1512 => x"33b3e700",
        1513 => x"33081841",
        1514 => x"33086840",
        1515 => x"33082803",
        1516 => x"33035703",
        1517 => x"b3382703",
        1518 => x"33086800",
        1519 => x"33072703",
        1520 => x"33081801",
        1521 => x"9358f841",
        1522 => x"93f83800",
        1523 => x"3387e800",
        1524 => x"b3381701",
        1525 => x"b3880801",
        1526 => x"9398e801",
        1527 => x"13572700",
        1528 => x"33e7e800",
        1529 => x"13184700",
        1530 => x"3307e840",
        1531 => x"13172700",
        1532 => x"338de740",
        1533 => x"eff0cf82",
        1534 => x"83260101",
        1535 => x"13070500",
        1536 => x"13880c00",
        1537 => x"93070d00",
        1538 => x"13060c00",
        1539 => x"93054bfb",
        1540 => x"13058101",
        1541 => x"ef00c015",
        1542 => x"13058101",
        1543 => x"efe0df9f",
        1544 => x"e3980be4",
        1545 => x"6ff05fe6",
        1546 => x"03a5c187",
        1547 => x"67800000",
        1548 => x"130101ff",
        1549 => x"23248100",
        1550 => x"23261100",
        1551 => x"93070000",
        1552 => x"13040500",
        1553 => x"63880700",
        1554 => x"93050000",
        1555 => x"97000000",
        1556 => x"e7000000",
        1557 => x"b7370000",
        1558 => x"03a50712",
        1559 => x"83278502",
        1560 => x"63840700",
        1561 => x"e7800700",
        1562 => x"13050400",
        1563 => x"ef100035",
        1564 => x"130101ff",
        1565 => x"23248100",
        1566 => x"23229100",
        1567 => x"37340000",
        1568 => x"b7340000",
        1569 => x"93874412",
        1570 => x"13044412",
        1571 => x"3304f440",
        1572 => x"23202101",
        1573 => x"23261100",
        1574 => x"13542440",
        1575 => x"93844412",
        1576 => x"13090000",
        1577 => x"63108904",
        1578 => x"b7340000",
        1579 => x"37340000",
        1580 => x"93874412",
        1581 => x"13044412",
        1582 => x"3304f440",
        1583 => x"13542440",
        1584 => x"93844412",
        1585 => x"13090000",
        1586 => x"63188902",
        1587 => x"8320c100",
        1588 => x"03248100",
        1589 => x"83244100",
        1590 => x"03290100",
        1591 => x"13010101",
        1592 => x"67800000",
        1593 => x"83a70400",
        1594 => x"13091900",
        1595 => x"93844400",
        1596 => x"e7800700",
        1597 => x"6ff01ffb",
        1598 => x"83a70400",
        1599 => x"13091900",
        1600 => x"93844400",
        1601 => x"e7800700",
        1602 => x"6ff01ffc",
        1603 => x"130101f6",
        1604 => x"232af108",
        1605 => x"b7070080",
        1606 => x"93c7f7ff",
        1607 => x"232ef100",
        1608 => x"2328f100",
        1609 => x"b707ffff",
        1610 => x"2326d108",
        1611 => x"2324b100",
        1612 => x"232cb100",
        1613 => x"93878720",
        1614 => x"9306c108",
        1615 => x"93058100",
        1616 => x"232e1106",
        1617 => x"232af100",
        1618 => x"2328e108",
        1619 => x"232c0109",
        1620 => x"232e1109",
        1621 => x"2322d100",
        1622 => x"ef00c040",
        1623 => x"83278100",
        1624 => x"23800700",
        1625 => x"8320c107",
        1626 => x"1301010a",
        1627 => x"67800000",
        1628 => x"130101f6",
        1629 => x"232af108",
        1630 => x"b7070080",
        1631 => x"93c7f7ff",
        1632 => x"232ef100",
        1633 => x"2328f100",
        1634 => x"b707ffff",
        1635 => x"93878720",
        1636 => x"232af100",
        1637 => x"2324a100",
        1638 => x"232ca100",
        1639 => x"03a5c187",
        1640 => x"2324c108",
        1641 => x"2326d108",
        1642 => x"13860500",
        1643 => x"93068108",
        1644 => x"93058100",
        1645 => x"232e1106",
        1646 => x"2328e108",
        1647 => x"232c0109",
        1648 => x"232e1109",
        1649 => x"2322d100",
        1650 => x"ef00c039",
        1651 => x"83278100",
        1652 => x"23800700",
        1653 => x"8320c107",
        1654 => x"1301010a",
        1655 => x"67800000",
        1656 => x"13860500",
        1657 => x"93050500",
        1658 => x"03a5c187",
        1659 => x"6f004000",
        1660 => x"130101ff",
        1661 => x"23248100",
        1662 => x"23229100",
        1663 => x"13040500",
        1664 => x"13850500",
        1665 => x"93050600",
        1666 => x"23261100",
        1667 => x"23a20188",
        1668 => x"ef10c01d",
        1669 => x"9307f0ff",
        1670 => x"6318f500",
        1671 => x"83a74188",
        1672 => x"63840700",
        1673 => x"2320f400",
        1674 => x"8320c100",
        1675 => x"03248100",
        1676 => x"83244100",
        1677 => x"13010101",
        1678 => x"67800000",
        1679 => x"130101fe",
        1680 => x"23282101",
        1681 => x"03a98500",
        1682 => x"232c8100",
        1683 => x"23263101",
        1684 => x"23225101",
        1685 => x"23206101",
        1686 => x"232e1100",
        1687 => x"232a9100",
        1688 => x"23244101",
        1689 => x"83aa0500",
        1690 => x"13840500",
        1691 => x"130b0600",
        1692 => x"93890600",
        1693 => x"63ec2609",
        1694 => x"8397c500",
        1695 => x"13f70748",
        1696 => x"63040708",
        1697 => x"03274401",
        1698 => x"93043000",
        1699 => x"83a50501",
        1700 => x"b384e402",
        1701 => x"13072000",
        1702 => x"b38aba40",
        1703 => x"130a0500",
        1704 => x"b3c4e402",
        1705 => x"13871600",
        1706 => x"33075701",
        1707 => x"63f4e400",
        1708 => x"93040700",
        1709 => x"93f70740",
        1710 => x"6386070a",
        1711 => x"93850400",
        1712 => x"13050a00",
        1713 => x"ef001067",
        1714 => x"13090500",
        1715 => x"630c050a",
        1716 => x"83250401",
        1717 => x"13860a00",
        1718 => x"eff05f9d",
        1719 => x"8357c400",
        1720 => x"93f7f7b7",
        1721 => x"93e70708",
        1722 => x"2316f400",
        1723 => x"23282401",
        1724 => x"232a9400",
        1725 => x"33095901",
        1726 => x"b3845441",
        1727 => x"23202401",
        1728 => x"23249400",
        1729 => x"13890900",
        1730 => x"63f42901",
        1731 => x"13890900",
        1732 => x"03250400",
        1733 => x"13060900",
        1734 => x"93050b00",
        1735 => x"eff01f9d",
        1736 => x"83278400",
        1737 => x"13050000",
        1738 => x"b3872741",
        1739 => x"2324f400",
        1740 => x"83270400",
        1741 => x"b3872701",
        1742 => x"2320f400",
        1743 => x"8320c101",
        1744 => x"03248101",
        1745 => x"83244101",
        1746 => x"03290101",
        1747 => x"8329c100",
        1748 => x"032a8100",
        1749 => x"832a4100",
        1750 => x"032b0100",
        1751 => x"13010102",
        1752 => x"67800000",
        1753 => x"13860400",
        1754 => x"13050a00",
        1755 => x"ef001071",
        1756 => x"13090500",
        1757 => x"e31c05f6",
        1758 => x"83250401",
        1759 => x"13050a00",
        1760 => x"ef00d04b",
        1761 => x"9307c000",
        1762 => x"2320fa00",
        1763 => x"8357c400",
        1764 => x"1305f0ff",
        1765 => x"93e70704",
        1766 => x"2316f400",
        1767 => x"6ff01ffa",
        1768 => x"83278600",
        1769 => x"130101fd",
        1770 => x"232e3101",
        1771 => x"23286101",
        1772 => x"23261102",
        1773 => x"23248102",
        1774 => x"23229102",
        1775 => x"23202103",
        1776 => x"232c4101",
        1777 => x"232a5101",
        1778 => x"23267101",
        1779 => x"23248101",
        1780 => x"23229101",
        1781 => x"2320a101",
        1782 => x"032b0600",
        1783 => x"93090600",
        1784 => x"63940712",
        1785 => x"13050000",
        1786 => x"8320c102",
        1787 => x"03248102",
        1788 => x"23a20900",
        1789 => x"83244102",
        1790 => x"03290102",
        1791 => x"8329c101",
        1792 => x"032a8101",
        1793 => x"832a4101",
        1794 => x"032b0101",
        1795 => x"832bc100",
        1796 => x"032c8100",
        1797 => x"832c4100",
        1798 => x"032d0100",
        1799 => x"13010103",
        1800 => x"67800000",
        1801 => x"832b0b00",
        1802 => x"032d4b00",
        1803 => x"130b8b00",
        1804 => x"03298400",
        1805 => x"832a0400",
        1806 => x"e3060dfe",
        1807 => x"63642d09",
        1808 => x"8317c400",
        1809 => x"13f70748",
        1810 => x"630e0706",
        1811 => x"83244401",
        1812 => x"83250401",
        1813 => x"b3049c02",
        1814 => x"b38aba40",
        1815 => x"13871a00",
        1816 => x"3307a701",
        1817 => x"b3c49403",
        1818 => x"63f4e400",
        1819 => x"93040700",
        1820 => x"93f70740",
        1821 => x"6388070a",
        1822 => x"93850400",
        1823 => x"13050a00",
        1824 => x"ef00504b",
        1825 => x"13090500",
        1826 => x"630e050a",
        1827 => x"83250401",
        1828 => x"13860a00",
        1829 => x"eff09f81",
        1830 => x"8357c400",
        1831 => x"93f7f7b7",
        1832 => x"93e70708",
        1833 => x"2316f400",
        1834 => x"23282401",
        1835 => x"232a9400",
        1836 => x"33095901",
        1837 => x"b3845441",
        1838 => x"23202401",
        1839 => x"23249400",
        1840 => x"13090d00",
        1841 => x"63742d01",
        1842 => x"13090d00",
        1843 => x"03250400",
        1844 => x"13060900",
        1845 => x"93850b00",
        1846 => x"eff05f81",
        1847 => x"83278400",
        1848 => x"b3872741",
        1849 => x"2324f400",
        1850 => x"83270400",
        1851 => x"b3872701",
        1852 => x"2320f400",
        1853 => x"83a78900",
        1854 => x"b387a741",
        1855 => x"23a4f900",
        1856 => x"e39207f2",
        1857 => x"6ff01fee",
        1858 => x"130a0500",
        1859 => x"13840500",
        1860 => x"930b0000",
        1861 => x"130d0000",
        1862 => x"130c3000",
        1863 => x"930c2000",
        1864 => x"6ff01ff1",
        1865 => x"13860400",
        1866 => x"13050a00",
        1867 => x"ef001055",
        1868 => x"13090500",
        1869 => x"e31a05f6",
        1870 => x"83250401",
        1871 => x"13050a00",
        1872 => x"ef00d02f",
        1873 => x"9307c000",
        1874 => x"2320fa00",
        1875 => x"8357c400",
        1876 => x"1305f0ff",
        1877 => x"93e70704",
        1878 => x"2316f400",
        1879 => x"23a40900",
        1880 => x"6ff09fe8",
        1881 => x"83d7c500",
        1882 => x"130101f5",
        1883 => x"2324810a",
        1884 => x"2322910a",
        1885 => x"2320210b",
        1886 => x"232c4109",
        1887 => x"2326110a",
        1888 => x"232e3109",
        1889 => x"232a5109",
        1890 => x"23286109",
        1891 => x"23267109",
        1892 => x"23248109",
        1893 => x"23229109",
        1894 => x"2320a109",
        1895 => x"232eb107",
        1896 => x"93f70708",
        1897 => x"130a0500",
        1898 => x"13890500",
        1899 => x"93040600",
        1900 => x"13840600",
        1901 => x"63880706",
        1902 => x"83a70501",
        1903 => x"63940706",
        1904 => x"93050004",
        1905 => x"ef001037",
        1906 => x"2320a900",
        1907 => x"2328a900",
        1908 => x"63160504",
        1909 => x"9307c000",
        1910 => x"2320fa00",
        1911 => x"1305f0ff",
        1912 => x"8320c10a",
        1913 => x"0324810a",
        1914 => x"8324410a",
        1915 => x"0329010a",
        1916 => x"8329c109",
        1917 => x"032a8109",
        1918 => x"832a4109",
        1919 => x"032b0109",
        1920 => x"832bc108",
        1921 => x"032c8108",
        1922 => x"832c4108",
        1923 => x"032d0108",
        1924 => x"832dc107",
        1925 => x"1301010b",
        1926 => x"67800000",
        1927 => x"93070004",
        1928 => x"232af900",
        1929 => x"93070002",
        1930 => x"a304f102",
        1931 => x"93070003",
        1932 => x"23220102",
        1933 => x"2305f102",
        1934 => x"23268100",
        1935 => x"930c5002",
        1936 => x"373b0000",
        1937 => x"b73b0000",
        1938 => x"373d0000",
        1939 => x"372c0000",
        1940 => x"930a0000",
        1941 => x"13840400",
        1942 => x"83470400",
        1943 => x"63840700",
        1944 => x"639c970d",
        1945 => x"b30d9440",
        1946 => x"63069402",
        1947 => x"93860d00",
        1948 => x"13860400",
        1949 => x"93050900",
        1950 => x"13050a00",
        1951 => x"eff01fbc",
        1952 => x"9307f0ff",
        1953 => x"6304f524",
        1954 => x"83274102",
        1955 => x"b387b701",
        1956 => x"2322f102",
        1957 => x"83470400",
        1958 => x"638a0722",
        1959 => x"9307f0ff",
        1960 => x"93041400",
        1961 => x"23280100",
        1962 => x"232e0100",
        1963 => x"232af100",
        1964 => x"232c0100",
        1965 => x"a3090104",
        1966 => x"23240106",
        1967 => x"930d1000",
        1968 => x"83c50400",
        1969 => x"13065000",
        1970 => x"1305cb08",
        1971 => x"ef00d014",
        1972 => x"83270101",
        1973 => x"13841400",
        1974 => x"63140506",
        1975 => x"13f70701",
        1976 => x"63060700",
        1977 => x"13070002",
        1978 => x"a309e104",
        1979 => x"13f78700",
        1980 => x"63060700",
        1981 => x"1307b002",
        1982 => x"a309e104",
        1983 => x"83c60400",
        1984 => x"1307a002",
        1985 => x"638ce604",
        1986 => x"8327c101",
        1987 => x"13840400",
        1988 => x"93060000",
        1989 => x"13069000",
        1990 => x"1305a000",
        1991 => x"03470400",
        1992 => x"93051400",
        1993 => x"130707fd",
        1994 => x"637ee608",
        1995 => x"63840604",
        1996 => x"232ef100",
        1997 => x"6f000004",
        1998 => x"13041400",
        1999 => x"6ff0dff1",
        2000 => x"1307cb08",
        2001 => x"3305e540",
        2002 => x"3395ad00",
        2003 => x"b3e7a700",
        2004 => x"2328f100",
        2005 => x"93040400",
        2006 => x"6ff09ff6",
        2007 => x"0327c100",
        2008 => x"93064700",
        2009 => x"03270700",
        2010 => x"2326d100",
        2011 => x"63420704",
        2012 => x"232ee100",
        2013 => x"03470400",
        2014 => x"9307e002",
        2015 => x"6314f708",
        2016 => x"03471400",
        2017 => x"9307a002",
        2018 => x"6318f704",
        2019 => x"8327c100",
        2020 => x"13042400",
        2021 => x"13874700",
        2022 => x"83a70700",
        2023 => x"2326e100",
        2024 => x"63d40700",
        2025 => x"9307f0ff",
        2026 => x"232af100",
        2027 => x"6f008005",
        2028 => x"3307e040",
        2029 => x"93e72700",
        2030 => x"232ee100",
        2031 => x"2328f100",
        2032 => x"6ff05ffb",
        2033 => x"b387a702",
        2034 => x"13840500",
        2035 => x"93061000",
        2036 => x"b387e700",
        2037 => x"6ff09ff4",
        2038 => x"13041400",
        2039 => x"232a0100",
        2040 => x"93060000",
        2041 => x"93070000",
        2042 => x"13069000",
        2043 => x"1305a000",
        2044 => x"03470400",
        2045 => x"93051400",
        2046 => x"130707fd",
        2047 => x"6372e608",
        2048 => x"e39406fa",
        2049 => x"83450400",
        2050 => x"13063000",
        2051 => x"13854b09",
        2052 => x"ef009000",
        2053 => x"63020502",
        2054 => x"93874b09",
        2055 => x"3305f540",
        2056 => x"83270101",
        2057 => x"13070004",
        2058 => x"3317a700",
        2059 => x"b3e7e700",
        2060 => x"13041400",
        2061 => x"2328f100",
        2062 => x"83450400",
        2063 => x"13066000",
        2064 => x"13058d09",
        2065 => x"93041400",
        2066 => x"2304b102",
        2067 => x"ef00c07c",
        2068 => x"63080508",
        2069 => x"63980a04",
        2070 => x"03270101",
        2071 => x"8327c100",
        2072 => x"13770710",
        2073 => x"63080702",
        2074 => x"93874700",
        2075 => x"2326f100",
        2076 => x"83274102",
        2077 => x"b3873701",
        2078 => x"2322f102",
        2079 => x"6ff09fdd",
        2080 => x"b387a702",
        2081 => x"13840500",
        2082 => x"93061000",
        2083 => x"b387e700",
        2084 => x"6ff01ff6",
        2085 => x"93877700",
        2086 => x"93f787ff",
        2087 => x"93878700",
        2088 => x"6ff0dffc",
        2089 => x"1307c100",
        2090 => x"9306cca3",
        2091 => x"13060900",
        2092 => x"93050101",
        2093 => x"13050a00",
        2094 => x"97000000",
        2095 => x"e7000000",
        2096 => x"9307f0ff",
        2097 => x"93090500",
        2098 => x"e314f5fa",
        2099 => x"8357c900",
        2100 => x"93f70704",
        2101 => x"e39407d0",
        2102 => x"03254102",
        2103 => x"6ff05fd0",
        2104 => x"1307c100",
        2105 => x"9306cca3",
        2106 => x"13060900",
        2107 => x"93050101",
        2108 => x"13050a00",
        2109 => x"ef00801b",
        2110 => x"6ff09ffc",
        2111 => x"130101fd",
        2112 => x"232a5101",
        2113 => x"83a70501",
        2114 => x"930a0700",
        2115 => x"03a78500",
        2116 => x"23248102",
        2117 => x"23202103",
        2118 => x"232e3101",
        2119 => x"232c4101",
        2120 => x"23261102",
        2121 => x"23229102",
        2122 => x"23286101",
        2123 => x"23267101",
        2124 => x"93090500",
        2125 => x"13840500",
        2126 => x"13090600",
        2127 => x"138a0600",
        2128 => x"63d4e700",
        2129 => x"93070700",
        2130 => x"2320f900",
        2131 => x"03473404",
        2132 => x"63060700",
        2133 => x"93871700",
        2134 => x"2320f900",
        2135 => x"83270400",
        2136 => x"93f70702",
        2137 => x"63880700",
        2138 => x"83270900",
        2139 => x"93872700",
        2140 => x"2320f900",
        2141 => x"83240400",
        2142 => x"93f46400",
        2143 => x"639e0400",
        2144 => x"130b9401",
        2145 => x"930bf0ff",
        2146 => x"8327c400",
        2147 => x"03270900",
        2148 => x"b387e740",
        2149 => x"63c2f408",
        2150 => x"83473404",
        2151 => x"b336f000",
        2152 => x"83270400",
        2153 => x"93f70702",
        2154 => x"6390070c",
        2155 => x"13063404",
        2156 => x"93050a00",
        2157 => x"13850900",
        2158 => x"e7800a00",
        2159 => x"9307f0ff",
        2160 => x"6308f506",
        2161 => x"83270400",
        2162 => x"13074000",
        2163 => x"93040000",
        2164 => x"93f76700",
        2165 => x"639ce700",
        2166 => x"8324c400",
        2167 => x"83270900",
        2168 => x"b384f440",
        2169 => x"63d40400",
        2170 => x"93040000",
        2171 => x"83278400",
        2172 => x"03270401",
        2173 => x"6356f700",
        2174 => x"b387e740",
        2175 => x"b384f400",
        2176 => x"13090000",
        2177 => x"1304a401",
        2178 => x"130bf0ff",
        2179 => x"63902409",
        2180 => x"13050000",
        2181 => x"6f000002",
        2182 => x"93061000",
        2183 => x"13060b00",
        2184 => x"93050a00",
        2185 => x"13850900",
        2186 => x"e7800a00",
        2187 => x"631a7503",
        2188 => x"1305f0ff",
        2189 => x"8320c102",
        2190 => x"03248102",
        2191 => x"83244102",
        2192 => x"03290102",
        2193 => x"8329c101",
        2194 => x"032a8101",
        2195 => x"832a4101",
        2196 => x"032b0101",
        2197 => x"832bc100",
        2198 => x"13010103",
        2199 => x"67800000",
        2200 => x"93841400",
        2201 => x"6ff05ff2",
        2202 => x"3307d400",
        2203 => x"13060003",
        2204 => x"a301c704",
        2205 => x"03475404",
        2206 => x"93871600",
        2207 => x"b307f400",
        2208 => x"93862600",
        2209 => x"a381e704",
        2210 => x"6ff05ff2",
        2211 => x"93061000",
        2212 => x"13060400",
        2213 => x"93050a00",
        2214 => x"13850900",
        2215 => x"e7800a00",
        2216 => x"e30865f9",
        2217 => x"13091900",
        2218 => x"6ff05ff6",
        2219 => x"130101fd",
        2220 => x"23248102",
        2221 => x"23229102",
        2222 => x"23202103",
        2223 => x"232e3101",
        2224 => x"23261102",
        2225 => x"232c4101",
        2226 => x"232a5101",
        2227 => x"23286101",
        2228 => x"83c88501",
        2229 => x"93078007",
        2230 => x"93040500",
        2231 => x"13840500",
        2232 => x"13090600",
        2233 => x"93890600",
        2234 => x"63ee1701",
        2235 => x"93072006",
        2236 => x"93863504",
        2237 => x"63ee1701",
        2238 => x"638a082a",
        2239 => x"93078005",
        2240 => x"638af820",
        2241 => x"930a2404",
        2242 => x"23011405",
        2243 => x"6f004004",
        2244 => x"9387d8f9",
        2245 => x"93f7f70f",
        2246 => x"13065001",
        2247 => x"e364f6fe",
        2248 => x"37360000",
        2249 => x"93972700",
        2250 => x"1306860c",
        2251 => x"b387c700",
        2252 => x"83a70700",
        2253 => x"67800700",
        2254 => x"83270700",
        2255 => x"938a2504",
        2256 => x"93864700",
        2257 => x"83a70700",
        2258 => x"2320d700",
        2259 => x"2381f504",
        2260 => x"93071000",
        2261 => x"6f004029",
        2262 => x"03a60500",
        2263 => x"83270700",
        2264 => x"13750608",
        2265 => x"93854700",
        2266 => x"630e0504",
        2267 => x"83a70700",
        2268 => x"2320b700",
        2269 => x"37370000",
        2270 => x"83254400",
        2271 => x"1308070a",
        2272 => x"63d2071e",
        2273 => x"1307d002",
        2274 => x"a301e404",
        2275 => x"2324b400",
        2276 => x"63d80504",
        2277 => x"b307f040",
        2278 => x"1307a000",
        2279 => x"938a0600",
        2280 => x"33f6e702",
        2281 => x"938afaff",
        2282 => x"3306c800",
        2283 => x"03460600",
        2284 => x"2380ca00",
        2285 => x"13860700",
        2286 => x"b3d7e702",
        2287 => x"e372e6fe",
        2288 => x"6f008009",
        2289 => x"83a70700",
        2290 => x"13750604",
        2291 => x"2320b700",
        2292 => x"e30205fa",
        2293 => x"93970701",
        2294 => x"93d70741",
        2295 => x"6ff09ff9",
        2296 => x"1376b6ff",
        2297 => x"2320c400",
        2298 => x"6ff0dffa",
        2299 => x"03a60500",
        2300 => x"83270700",
        2301 => x"13750608",
        2302 => x"93854700",
        2303 => x"63080500",
        2304 => x"2320b700",
        2305 => x"83a70700",
        2306 => x"6f004001",
        2307 => x"13760604",
        2308 => x"2320b700",
        2309 => x"e30806fe",
        2310 => x"83d70700",
        2311 => x"37380000",
        2312 => x"1307f006",
        2313 => x"1308080a",
        2314 => x"639ae812",
        2315 => x"13078000",
        2316 => x"a3010404",
        2317 => x"03264400",
        2318 => x"2324c400",
        2319 => x"e34006f6",
        2320 => x"83250400",
        2321 => x"93f5b5ff",
        2322 => x"2320b400",
        2323 => x"e39807f4",
        2324 => x"938a0600",
        2325 => x"e31406f4",
        2326 => x"93078000",
        2327 => x"6314f702",
        2328 => x"83270400",
        2329 => x"93f71700",
        2330 => x"638e0700",
        2331 => x"03274400",
        2332 => x"83270401",
        2333 => x"63c8e700",
        2334 => x"93070003",
        2335 => x"a38ffafe",
        2336 => x"938afaff",
        2337 => x"b3865641",
        2338 => x"2328d400",
        2339 => x"13870900",
        2340 => x"93060900",
        2341 => x"1306c100",
        2342 => x"93050400",
        2343 => x"13850400",
        2344 => x"eff0dfc5",
        2345 => x"130af0ff",
        2346 => x"63164515",
        2347 => x"1305f0ff",
        2348 => x"8320c102",
        2349 => x"03248102",
        2350 => x"83244102",
        2351 => x"03290102",
        2352 => x"8329c101",
        2353 => x"032a8101",
        2354 => x"832a4101",
        2355 => x"032b0101",
        2356 => x"13010103",
        2357 => x"67800000",
        2358 => x"83a70500",
        2359 => x"93e70702",
        2360 => x"23a0f500",
        2361 => x"37380000",
        2362 => x"93088007",
        2363 => x"1308480b",
        2364 => x"03260400",
        2365 => x"a3021405",
        2366 => x"83270700",
        2367 => x"13750608",
        2368 => x"93854700",
        2369 => x"630e0500",
        2370 => x"2320b700",
        2371 => x"83a70700",
        2372 => x"6f000002",
        2373 => x"37380000",
        2374 => x"1308080a",
        2375 => x"6ff05ffd",
        2376 => x"13750604",
        2377 => x"2320b700",
        2378 => x"e30205fe",
        2379 => x"83d70700",
        2380 => x"13771600",
        2381 => x"63060700",
        2382 => x"13660602",
        2383 => x"2320c400",
        2384 => x"63860700",
        2385 => x"13070001",
        2386 => x"6ff09fee",
        2387 => x"03270400",
        2388 => x"1377f7fd",
        2389 => x"2320e400",
        2390 => x"6ff0dffe",
        2391 => x"1307a000",
        2392 => x"6ff01fed",
        2393 => x"1308070a",
        2394 => x"1307a000",
        2395 => x"6ff09fec",
        2396 => x"03a60500",
        2397 => x"83270700",
        2398 => x"83a54501",
        2399 => x"13780608",
        2400 => x"13854700",
        2401 => x"630a0800",
        2402 => x"2320a700",
        2403 => x"83a70700",
        2404 => x"23a0b700",
        2405 => x"6f008001",
        2406 => x"2320a700",
        2407 => x"13760604",
        2408 => x"83a70700",
        2409 => x"e30606fe",
        2410 => x"2390b700",
        2411 => x"23280400",
        2412 => x"938a0600",
        2413 => x"6ff09fed",
        2414 => x"83270700",
        2415 => x"03a64500",
        2416 => x"93050000",
        2417 => x"93864700",
        2418 => x"2320d700",
        2419 => x"83aa0700",
        2420 => x"13850a00",
        2421 => x"ef004024",
        2422 => x"63060500",
        2423 => x"33055541",
        2424 => x"2322a400",
        2425 => x"83274400",
        2426 => x"2328f400",
        2427 => x"a3010404",
        2428 => x"6ff0dfe9",
        2429 => x"83260401",
        2430 => x"13860a00",
        2431 => x"93050900",
        2432 => x"13850400",
        2433 => x"e7800900",
        2434 => x"e30245eb",
        2435 => x"83270400",
        2436 => x"93f72700",
        2437 => x"63940704",
        2438 => x"8327c100",
        2439 => x"0325c400",
        2440 => x"e358f5e8",
        2441 => x"13850700",
        2442 => x"6ff09fe8",
        2443 => x"93061000",
        2444 => x"13860a00",
        2445 => x"93050900",
        2446 => x"13850400",
        2447 => x"e7800900",
        2448 => x"e30665e7",
        2449 => x"130a1a00",
        2450 => x"8327c400",
        2451 => x"0327c100",
        2452 => x"b387e740",
        2453 => x"e34cfafc",
        2454 => x"6ff01ffc",
        2455 => x"130a0000",
        2456 => x"930a9401",
        2457 => x"130bf0ff",
        2458 => x"6ff01ffe",
        2459 => x"130101ff",
        2460 => x"23248100",
        2461 => x"13840500",
        2462 => x"83a50500",
        2463 => x"23229100",
        2464 => x"23261100",
        2465 => x"93040500",
        2466 => x"63840500",
        2467 => x"eff01ffe",
        2468 => x"93050400",
        2469 => x"03248100",
        2470 => x"8320c100",
        2471 => x"13850400",
        2472 => x"83244100",
        2473 => x"13010101",
        2474 => x"6f004019",
        2475 => x"83a7c187",
        2476 => x"6382a716",
        2477 => x"83274502",
        2478 => x"130101fe",
        2479 => x"232c8100",
        2480 => x"232e1100",
        2481 => x"232a9100",
        2482 => x"23282101",
        2483 => x"23263101",
        2484 => x"13040500",
        2485 => x"638a0704",
        2486 => x"83a7c700",
        2487 => x"638c0702",
        2488 => x"93040000",
        2489 => x"13090008",
        2490 => x"83274402",
        2491 => x"83a7c700",
        2492 => x"b3879700",
        2493 => x"83a50700",
        2494 => x"6396050e",
        2495 => x"93844400",
        2496 => x"e39424ff",
        2497 => x"83274402",
        2498 => x"13050400",
        2499 => x"83a5c700",
        2500 => x"ef00c012",
        2501 => x"83274402",
        2502 => x"83a50700",
        2503 => x"63860500",
        2504 => x"13050400",
        2505 => x"ef008011",
        2506 => x"83254401",
        2507 => x"63860500",
        2508 => x"13050400",
        2509 => x"ef008010",
        2510 => x"83254402",
        2511 => x"63860500",
        2512 => x"13050400",
        2513 => x"ef00800f",
        2514 => x"83258403",
        2515 => x"63860500",
        2516 => x"13050400",
        2517 => x"ef00800e",
        2518 => x"8325c403",
        2519 => x"63860500",
        2520 => x"13050400",
        2521 => x"ef00800d",
        2522 => x"83250404",
        2523 => x"63860500",
        2524 => x"13050400",
        2525 => x"ef00800c",
        2526 => x"8325c405",
        2527 => x"63860500",
        2528 => x"13050400",
        2529 => x"ef00800b",
        2530 => x"83258405",
        2531 => x"63860500",
        2532 => x"13050400",
        2533 => x"ef00800a",
        2534 => x"83254403",
        2535 => x"63860500",
        2536 => x"13050400",
        2537 => x"ef008009",
        2538 => x"83278401",
        2539 => x"63860704",
        2540 => x"83278402",
        2541 => x"13050400",
        2542 => x"e7800700",
        2543 => x"83258404",
        2544 => x"638c0502",
        2545 => x"13050400",
        2546 => x"03248101",
        2547 => x"8320c101",
        2548 => x"83244101",
        2549 => x"03290101",
        2550 => x"8329c100",
        2551 => x"13010102",
        2552 => x"6ff0dfe8",
        2553 => x"83a90500",
        2554 => x"13050400",
        2555 => x"ef000005",
        2556 => x"93850900",
        2557 => x"6ff05ff0",
        2558 => x"8320c101",
        2559 => x"03248101",
        2560 => x"83244101",
        2561 => x"03290101",
        2562 => x"8329c100",
        2563 => x"13010102",
        2564 => x"67800000",
        2565 => x"67800000",
        2566 => x"93f5f50f",
        2567 => x"3306c500",
        2568 => x"6316c500",
        2569 => x"13050000",
        2570 => x"67800000",
        2571 => x"83470500",
        2572 => x"e38cb7fe",
        2573 => x"13051500",
        2574 => x"6ff09ffe",
        2575 => x"638a050e",
        2576 => x"83a7c5ff",
        2577 => x"130101fe",
        2578 => x"232c8100",
        2579 => x"232e1100",
        2580 => x"1384c5ff",
        2581 => x"63d40700",
        2582 => x"3304f400",
        2583 => x"2326a100",
        2584 => x"ef008033",
        2585 => x"83a7c188",
        2586 => x"0325c100",
        2587 => x"639e0700",
        2588 => x"23220400",
        2589 => x"23a68188",
        2590 => x"03248101",
        2591 => x"8320c101",
        2592 => x"13010102",
        2593 => x"6f008031",
        2594 => x"6374f402",
        2595 => x"03260400",
        2596 => x"b306c400",
        2597 => x"639ad700",
        2598 => x"83a60700",
        2599 => x"83a74700",
        2600 => x"b386c600",
        2601 => x"2320d400",
        2602 => x"2322f400",
        2603 => x"6ff09ffc",
        2604 => x"13870700",
        2605 => x"83a74700",
        2606 => x"63840700",
        2607 => x"e37af4fe",
        2608 => x"83260700",
        2609 => x"3306d700",
        2610 => x"63188602",
        2611 => x"03260400",
        2612 => x"b386c600",
        2613 => x"2320d700",
        2614 => x"3306d700",
        2615 => x"e39ec7f8",
        2616 => x"03a60700",
        2617 => x"83a74700",
        2618 => x"b306d600",
        2619 => x"2320d700",
        2620 => x"2322f700",
        2621 => x"6ff05ff8",
        2622 => x"6378c400",
        2623 => x"9307c000",
        2624 => x"2320f500",
        2625 => x"6ff05ff7",
        2626 => x"03260400",
        2627 => x"b306c400",
        2628 => x"639ad700",
        2629 => x"83a60700",
        2630 => x"83a74700",
        2631 => x"b386c600",
        2632 => x"2320d400",
        2633 => x"2322f400",
        2634 => x"23228700",
        2635 => x"6ff0dff4",
        2636 => x"67800000",
        2637 => x"130101fe",
        2638 => x"232a9100",
        2639 => x"93843500",
        2640 => x"93f4c4ff",
        2641 => x"23282101",
        2642 => x"232e1100",
        2643 => x"232c8100",
        2644 => x"23263101",
        2645 => x"93848400",
        2646 => x"9307c000",
        2647 => x"13090500",
        2648 => x"63f0f406",
        2649 => x"9304c000",
        2650 => x"63eeb404",
        2651 => x"13050900",
        2652 => x"ef008022",
        2653 => x"03a7c188",
        2654 => x"13040700",
        2655 => x"63180406",
        2656 => x"83a78188",
        2657 => x"639a0700",
        2658 => x"93050000",
        2659 => x"13050900",
        2660 => x"ef00001c",
        2661 => x"23a4a188",
        2662 => x"93850400",
        2663 => x"13050900",
        2664 => x"ef00001b",
        2665 => x"9309f0ff",
        2666 => x"631a350b",
        2667 => x"9307c000",
        2668 => x"2320f900",
        2669 => x"13050900",
        2670 => x"ef00401e",
        2671 => x"6f000001",
        2672 => x"e3d404fa",
        2673 => x"9307c000",
        2674 => x"2320f900",
        2675 => x"13050000",
        2676 => x"8320c101",
        2677 => x"03248101",
        2678 => x"83244101",
        2679 => x"03290101",
        2680 => x"8329c100",
        2681 => x"13010102",
        2682 => x"67800000",
        2683 => x"83270400",
        2684 => x"b3879740",
        2685 => x"63ce0704",
        2686 => x"1306b000",
        2687 => x"637af600",
        2688 => x"2320f400",
        2689 => x"3304f400",
        2690 => x"23209400",
        2691 => x"6f000001",
        2692 => x"83274400",
        2693 => x"631a8702",
        2694 => x"23a6f188",
        2695 => x"13050900",
        2696 => x"ef00c017",
        2697 => x"1305b400",
        2698 => x"93074400",
        2699 => x"137585ff",
        2700 => x"3307f540",
        2701 => x"e30ef5f8",
        2702 => x"3304e400",
        2703 => x"b387a740",
        2704 => x"2320f400",
        2705 => x"6ff0dff8",
        2706 => x"2322f700",
        2707 => x"6ff01ffd",
        2708 => x"13070400",
        2709 => x"03244400",
        2710 => x"6ff05ff2",
        2711 => x"13043500",
        2712 => x"1374c4ff",
        2713 => x"e30285fa",
        2714 => x"b305a440",
        2715 => x"13050900",
        2716 => x"ef00000e",
        2717 => x"e31a35f9",
        2718 => x"6ff05ff3",
        2719 => x"130101fe",
        2720 => x"232c8100",
        2721 => x"232e1100",
        2722 => x"232a9100",
        2723 => x"23282101",
        2724 => x"23263101",
        2725 => x"23244101",
        2726 => x"13040600",
        2727 => x"63940502",
        2728 => x"03248101",
        2729 => x"8320c101",
        2730 => x"83244101",
        2731 => x"03290101",
        2732 => x"8329c100",
        2733 => x"032a8100",
        2734 => x"93050600",
        2735 => x"13010102",
        2736 => x"6ff05fe7",
        2737 => x"63180602",
        2738 => x"eff05fd7",
        2739 => x"93040000",
        2740 => x"8320c101",
        2741 => x"03248101",
        2742 => x"03290101",
        2743 => x"8329c100",
        2744 => x"032a8100",
        2745 => x"13850400",
        2746 => x"83244101",
        2747 => x"13010102",
        2748 => x"67800000",
        2749 => x"130a0500",
        2750 => x"93840500",
        2751 => x"ef00400a",
        2752 => x"13090500",
        2753 => x"63668500",
        2754 => x"93571500",
        2755 => x"e3e287fc",
        2756 => x"93050400",
        2757 => x"13050a00",
        2758 => x"eff0dfe1",
        2759 => x"93090500",
        2760 => x"e30605fa",
        2761 => x"13060400",
        2762 => x"63748900",
        2763 => x"13060900",
        2764 => x"93850400",
        2765 => x"13850900",
        2766 => x"efe05f97",
        2767 => x"93850400",
        2768 => x"13050a00",
        2769 => x"eff09fcf",
        2770 => x"93840900",
        2771 => x"6ff05ff8",
        2772 => x"130101ff",
        2773 => x"23248100",
        2774 => x"23229100",
        2775 => x"13040500",
        2776 => x"13850500",
        2777 => x"23261100",
        2778 => x"23a20188",
        2779 => x"ef00000c",
        2780 => x"9307f0ff",
        2781 => x"6318f500",
        2782 => x"83a74188",
        2783 => x"63840700",
        2784 => x"2320f400",
        2785 => x"8320c100",
        2786 => x"03248100",
        2787 => x"83244100",
        2788 => x"13010101",
        2789 => x"67800000",
        2790 => x"67800000",
        2791 => x"67800000",
        2792 => x"83a7c5ff",
        2793 => x"1385c7ff",
        2794 => x"63d80700",
        2795 => x"b385a500",
        2796 => x"83a70500",
        2797 => x"3305f500",
        2798 => x"67800000",
        2799 => x"9308d005",
        2800 => x"73000000",
        2801 => x"63520502",
        2802 => x"130101ff",
        2803 => x"23248100",
        2804 => x"13040500",
        2805 => x"23261100",
        2806 => x"33048040",
        2807 => x"efe0dfc4",
        2808 => x"23208500",
        2809 => x"6f000000",
        2810 => x"6f000000",
        2811 => x"130101ff",
        2812 => x"23261100",
        2813 => x"23248100",
        2814 => x"9308900a",
        2815 => x"73000000",
        2816 => x"13040500",
        2817 => x"635a0500",
        2818 => x"33048040",
        2819 => x"efe0dfc1",
        2820 => x"23208500",
        2821 => x"1304f0ff",
        2822 => x"8320c100",
        2823 => x"13050400",
        2824 => x"03248100",
        2825 => x"13010101",
        2826 => x"67800000",
        2827 => x"03a70189",
        2828 => x"130101ff",
        2829 => x"23261100",
        2830 => x"93070500",
        2831 => x"631c0702",
        2832 => x"9308600d",
        2833 => x"13050000",
        2834 => x"73000000",
        2835 => x"1307f0ff",
        2836 => x"6310e502",
        2837 => x"efe05fbd",
        2838 => x"9307c000",
        2839 => x"2320f500",
        2840 => x"1305f0ff",
        2841 => x"8320c100",
        2842 => x"13010101",
        2843 => x"67800000",
        2844 => x"23a8a188",
        2845 => x"03a70189",
        2846 => x"9308600d",
        2847 => x"b387e700",
        2848 => x"13850700",
        2849 => x"73000000",
        2850 => x"e316f5fc",
        2851 => x"23a8a188",
        2852 => x"13050700",
        2853 => x"6ff01ffd",
        2854 => x"10000000",
        2855 => x"00000000",
        2856 => x"037a5200",
        2857 => x"017c0101",
        2858 => x"1b0d0200",
        2859 => x"10000000",
        2860 => x"18000000",
        2861 => x"6cdbffff",
        2862 => x"78040000",
        2863 => x"00000000",
        2864 => x"10000000",
        2865 => x"00000000",
        2866 => x"037a5200",
        2867 => x"017c0101",
        2868 => x"1b0d0200",
        2869 => x"10000000",
        2870 => x"18000000",
        2871 => x"bcdfffff",
        2872 => x"30040000",
        2873 => x"00000000",
        2874 => x"10000000",
        2875 => x"00000000",
        2876 => x"037a5200",
        2877 => x"017c0101",
        2878 => x"1b0d0200",
        2879 => x"10000000",
        2880 => x"18000000",
        2881 => x"c4e3ffff",
        2882 => x"e4030000",
        2883 => x"00000000",
        2884 => x"a4030000",
        2885 => x"d4020000",
        2886 => x"d4020000",
        2887 => x"d4020000",
        2888 => x"d4020000",
        2889 => x"4c030000",
        2890 => x"d4020000",
        2891 => x"14030000",
        2892 => x"d4020000",
        2893 => x"d4020000",
        2894 => x"14030000",
        2895 => x"d4020000",
        2896 => x"d4020000",
        2897 => x"d4020000",
        2898 => x"d4020000",
        2899 => x"d4020000",
        2900 => x"d4020000",
        2901 => x"d4020000",
        2902 => x"74030000",
        2903 => x"10060000",
        2904 => x"ec050000",
        2905 => x"04060000",
        2906 => x"f8050000",
        2907 => x"40050000",
        2908 => x"40050000",
        2909 => x"40050000",
        2910 => x"54060000",
        2911 => x"40050000",
        2912 => x"40050000",
        2913 => x"40050000",
        2914 => x"40050000",
        2915 => x"40050000",
        2916 => x"40050000",
        2917 => x"40050000",
        2918 => x"1c060000",
        2919 => x"b8060000",
        2920 => x"70060000",
        2921 => x"70060000",
        2922 => x"70060000",
        2923 => x"70060000",
        2924 => x"ac060000",
        2925 => x"f8060000",
        2926 => x"d0060000",
        2927 => x"70060000",
        2928 => x"70060000",
        2929 => x"70060000",
        2930 => x"70060000",
        2931 => x"70060000",
        2932 => x"70060000",
        2933 => x"70060000",
        2934 => x"70060000",
        2935 => x"70060000",
        2936 => x"70060000",
        2937 => x"70060000",
        2938 => x"70060000",
        2939 => x"70060000",
        2940 => x"70060000",
        2941 => x"98060000",
        2942 => x"98060000",
        2943 => x"70060000",
        2944 => x"70060000",
        2945 => x"70060000",
        2946 => x"70060000",
        2947 => x"70060000",
        2948 => x"70060000",
        2949 => x"70060000",
        2950 => x"70060000",
        2951 => x"70060000",
        2952 => x"70060000",
        2953 => x"70060000",
        2954 => x"70060000",
        2955 => x"ac060000",
        2956 => x"b8060000",
        2957 => x"74070000",
        2958 => x"5c070000",
        2959 => x"70060000",
        2960 => x"70060000",
        2961 => x"70060000",
        2962 => x"70060000",
        2963 => x"70060000",
        2964 => x"70060000",
        2965 => x"44070000",
        2966 => x"70060000",
        2967 => x"70060000",
        2968 => x"70060000",
        2969 => x"70060000",
        2970 => x"98060000",
        2971 => x"98060000",
        2972 => x"00010202",
        2973 => x"03030303",
        2974 => x"04040404",
        2975 => x"04040404",
        2976 => x"05050505",
        2977 => x"05050505",
        2978 => x"05050505",
        2979 => x"05050505",
        2980 => x"06060606",
        2981 => x"06060606",
        2982 => x"06060606",
        2983 => x"06060606",
        2984 => x"06060606",
        2985 => x"06060606",
        2986 => x"06060606",
        2987 => x"06060606",
        2988 => x"07070707",
        2989 => x"07070707",
        2990 => x"07070707",
        2991 => x"07070707",
        2992 => x"07070707",
        2993 => x"07070707",
        2994 => x"07070707",
        2995 => x"07070707",
        2996 => x"07070707",
        2997 => x"07070707",
        2998 => x"07070707",
        2999 => x"07070707",
        3000 => x"07070707",
        3001 => x"07070707",
        3002 => x"07070707",
        3003 => x"07070707",
        3004 => x"08080808",
        3005 => x"08080808",
        3006 => x"08080808",
        3007 => x"08080808",
        3008 => x"08080808",
        3009 => x"08080808",
        3010 => x"08080808",
        3011 => x"08080808",
        3012 => x"08080808",
        3013 => x"08080808",
        3014 => x"08080808",
        3015 => x"08080808",
        3016 => x"08080808",
        3017 => x"08080808",
        3018 => x"08080808",
        3019 => x"08080808",
        3020 => x"08080808",
        3021 => x"08080808",
        3022 => x"08080808",
        3023 => x"08080808",
        3024 => x"08080808",
        3025 => x"08080808",
        3026 => x"08080808",
        3027 => x"08080808",
        3028 => x"08080808",
        3029 => x"08080808",
        3030 => x"08080808",
        3031 => x"08080808",
        3032 => x"08080808",
        3033 => x"08080808",
        3034 => x"08080808",
        3035 => x"08080808",
        3036 => x"0d0a4542",
        3037 => x"5245414b",
        3038 => x"21206d69",
        3039 => x"70203d20",
        3040 => x"00000000",
        3041 => x"0d0a0d0a",
        3042 => x"44697370",
        3043 => x"6c617969",
        3044 => x"6e672074",
        3045 => x"68652074",
        3046 => x"696d6520",
        3047 => x"70617373",
        3048 => x"65642073",
        3049 => x"696e6365",
        3050 => x"20726573",
        3051 => x"65740d0a",
        3052 => x"0d0a0000",
        3053 => x"2530356c",
        3054 => x"643a2530",
        3055 => x"366c6420",
        3056 => x"20202530",
        3057 => x"326c643a",
        3058 => x"2530326c",
        3059 => x"643a2530",
        3060 => x"326c640d",
        3061 => x"00000000",
        3062 => x"696e7465",
        3063 => x"72727570",
        3064 => x"745f6469",
        3065 => x"72656374",
        3066 => x"00000000",
        3067 => x"54485541",
        3068 => x"53205249",
        3069 => x"53432d56",
        3070 => x"20525633",
        3071 => x"32494d20",
        3072 => x"62617265",
        3073 => x"206d6574",
        3074 => x"616c2070",
        3075 => x"726f6365",
        3076 => x"73736f72",
        3077 => x"00000000",
        3078 => x"54686520",
        3079 => x"48616775",
        3080 => x"6520556e",
        3081 => x"69766572",
        3082 => x"73697479",
        3083 => x"206f6620",
        3084 => x"4170706c",
        3085 => x"69656420",
        3086 => x"53636965",
        3087 => x"6e636573",
        3088 => x"00000000",
        3089 => x"44657061",
        3090 => x"72746d65",
        3091 => x"6e74206f",
        3092 => x"6620456c",
        3093 => x"65637472",
        3094 => x"6963616c",
        3095 => x"20456e67",
        3096 => x"696e6565",
        3097 => x"72696e67",
        3098 => x"00000000",
        3099 => x"4a2e452e",
        3100 => x"4a2e206f",
        3101 => x"70206465",
        3102 => x"6e204272",
        3103 => x"6f757700",
        3104 => x"3c627265",
        3105 => x"616b3e0d",
        3106 => x"0a000000",
        3107 => x"232d302b",
        3108 => x"20000000",
        3109 => x"686c4c00",
        3110 => x"65666745",
        3111 => x"46470000",
        3112 => x"30313233",
        3113 => x"34353637",
        3114 => x"38394142",
        3115 => x"43444546",
        3116 => x"00000000",
        3117 => x"30313233",
        3118 => x"34353637",
        3119 => x"38396162",
        3120 => x"63646566",
        3121 => x"00000000",
        3122 => x"38230000",
        3123 => x"58230000",
        3124 => x"04230000",
        3125 => x"04230000",
        3126 => x"04230000",
        3127 => x"04230000",
        3128 => x"58230000",
        3129 => x"04230000",
        3130 => x"04230000",
        3131 => x"04230000",
        3132 => x"04230000",
        3133 => x"70250000",
        3134 => x"ec230000",
        3135 => x"d8240000",
        3136 => x"04230000",
        3137 => x"04230000",
        3138 => x"b8250000",
        3139 => x"04230000",
        3140 => x"ec230000",
        3141 => x"04230000",
        3142 => x"04230000",
        3143 => x"e4240000",
        3144 => x"18000020",
        3145 => x"d82f0000",
        3146 => x"ec2f0000",
        3147 => x"18300000",
        3148 => x"44300000",
        3149 => x"6c300000",
        3150 => x"00000000",
        3151 => x"00000000",
        3152 => x"00000000",
        3153 => x"00000000",
        3154 => x"00000000",
        3155 => x"00000000",
        3156 => x"00000000",
        3157 => x"00000000",
        3158 => x"00000000",
        3159 => x"00000000",
        3160 => x"00000000",
        3161 => x"00000000",
        3162 => x"00000000",
        3163 => x"00000000",
        3164 => x"00000000",
        3165 => x"00000000",
        3166 => x"00000000",
        3167 => x"00000000",
        3168 => x"00000000",
        3169 => x"00000000",
        3170 => x"00000000",
        3171 => x"00000000",
        3172 => x"00000000",
        3173 => x"00000000",
        3174 => x"00000000",
        3175 => x"80000020",
        3176 => x"18000020",
        others => (others => '0')
    );
end package processor_common_rom;
