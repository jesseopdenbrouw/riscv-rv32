-- srec2vhdl table generator
-- for input file interrupt_direct.srec

library ieee;
use ieee.std_logic_1164.all;

library work;
use work.processor_common.all;

package processor_common_rom is
    constant rom_contents : rom_type := (
           0 => x"97110020",
           1 => x"93810180",
           2 => x"17810020",
           3 => x"130181ff",
           4 => x"97020000",
           5 => x"9382421f",
           6 => x"73905230",
           7 => x"13860188",
           8 => x"93874189",
           9 => x"637af600",
          10 => x"3386c740",
          11 => x"93050000",
          12 => x"13850188",
          13 => x"ef10802d",
          14 => x"37050020",
          15 => x"13060500",
          16 => x"93870188",
          17 => x"637cf600",
          18 => x"b7350000",
          19 => x"3386c740",
          20 => x"938585f0",
          21 => x"13050500",
          22 => x"ef100029",
          23 => x"ef100065",
          24 => x"b7050020",
          25 => x"13060000",
          26 => x"93850500",
          27 => x"13055000",
          28 => x"ef10402f",
          29 => x"ef10805f",
          30 => x"6f008055",
          31 => x"130101ff",
          32 => x"23261100",
          33 => x"ef008057",
          34 => x"8320c100",
          35 => x"13051000",
          36 => x"13010101",
          37 => x"67800000",
          38 => x"37350000",
          39 => x"130101ff",
          40 => x"130505d6",
          41 => x"23261100",
          42 => x"23248100",
          43 => x"23229100",
          44 => x"23202101",
          45 => x"ef008056",
          46 => x"73294034",
          47 => x"93040002",
          48 => x"37040080",
          49 => x"33758900",
          50 => x"3335a000",
          51 => x"13050503",
          52 => x"9384f4ff",
          53 => x"ef008052",
          54 => x"13541400",
          55 => x"e39404fe",
          56 => x"03248100",
          57 => x"8320c100",
          58 => x"83244100",
          59 => x"03290100",
          60 => x"37350000",
          61 => x"130505da",
          62 => x"13010101",
          63 => x"6f000052",
          64 => x"b70700f0",
          65 => x"03a74708",
          66 => x"1377f7fe",
          67 => x"23a2e708",
          68 => x"03a74700",
          69 => x"13471700",
          70 => x"23a2e700",
          71 => x"67800000",
          72 => x"370700f0",
          73 => x"83274700",
          74 => x"93e70720",
          75 => x"2322f700",
          76 => x"6f000000",
          77 => x"b70700f0",
          78 => x"83a6470f",
          79 => x"03a6070f",
          80 => x"03a7470f",
          81 => x"e31ad7fe",
          82 => x"b7860100",
          83 => x"9305f0ff",
          84 => x"9386066a",
          85 => x"23aeb70e",
          86 => x"b306d600",
          87 => x"23acb70e",
          88 => x"33b6c600",
          89 => x"23acd70e",
          90 => x"3306e600",
          91 => x"23aec70e",
          92 => x"03a74700",
          93 => x"13472700",
          94 => x"23a2e700",
          95 => x"67800000",
          96 => x"370700f0",
          97 => x"8327c702",
          98 => x"93f74700",
          99 => x"638a0700",
         100 => x"83274700",
         101 => x"93c78700",
         102 => x"2322f700",
         103 => x"83270702",
         104 => x"67800000",
         105 => x"b70700f0",
         106 => x"03a7470a",
         107 => x"1377f7f0",
         108 => x"23a2e70a",
         109 => x"03a74700",
         110 => x"13474700",
         111 => x"23a2e700",
         112 => x"67800000",
         113 => x"b70700f0",
         114 => x"03a74706",
         115 => x"137777ff",
         116 => x"23a2e706",
         117 => x"03a74700",
         118 => x"13470701",
         119 => x"23a2e700",
         120 => x"67800000",
         121 => x"b70700f0",
         122 => x"03a74704",
         123 => x"137777fe",
         124 => x"23a2e704",
         125 => x"03a74700",
         126 => x"13470702",
         127 => x"23a2e700",
         128 => x"67800000",
         129 => x"6f000000",
         130 => x"13050000",
         131 => x"67800000",
         132 => x"13050000",
         133 => x"67800000",
         134 => x"130101f8",
         135 => x"23221100",
         136 => x"23242100",
         137 => x"23263100",
         138 => x"23284100",
         139 => x"232a5100",
         140 => x"232c6100",
         141 => x"232e7100",
         142 => x"23208102",
         143 => x"23229102",
         144 => x"2324a102",
         145 => x"2326b102",
         146 => x"2328c102",
         147 => x"232ad102",
         148 => x"232ce102",
         149 => x"232ef102",
         150 => x"23200105",
         151 => x"23221105",
         152 => x"23242105",
         153 => x"23263105",
         154 => x"23284105",
         155 => x"232a5105",
         156 => x"232c6105",
         157 => x"232e7105",
         158 => x"23208107",
         159 => x"23229107",
         160 => x"2324a107",
         161 => x"2326b107",
         162 => x"2328c107",
         163 => x"232ad107",
         164 => x"232ce107",
         165 => x"232ef107",
         166 => x"f3272034",
         167 => x"37070080",
         168 => x"93067700",
         169 => x"6386d70e",
         170 => x"9306b000",
         171 => x"63fef602",
         172 => x"9346f7fe",
         173 => x"b386d700",
         174 => x"13064000",
         175 => x"636ad602",
         176 => x"1347e7fe",
         177 => x"b387e700",
         178 => x"13073000",
         179 => x"6364f714",
         180 => x"37370000",
         181 => x"93972700",
         182 => x"1307c7b4",
         183 => x"b387e700",
         184 => x"83a70700",
         185 => x"67800700",
         186 => x"13071000",
         187 => x"6364f708",
         188 => x"03258102",
         189 => x"832fc107",
         190 => x"032f8107",
         191 => x"832e4107",
         192 => x"032e0107",
         193 => x"832dc106",
         194 => x"032d8106",
         195 => x"832c4106",
         196 => x"032c0106",
         197 => x"832bc105",
         198 => x"032b8105",
         199 => x"832a4105",
         200 => x"032a0105",
         201 => x"8329c104",
         202 => x"03298104",
         203 => x"83284104",
         204 => x"03280104",
         205 => x"8327c103",
         206 => x"03278103",
         207 => x"83264103",
         208 => x"03260103",
         209 => x"8325c102",
         210 => x"83244102",
         211 => x"03240102",
         212 => x"8323c101",
         213 => x"03238101",
         214 => x"83224101",
         215 => x"03220101",
         216 => x"8321c100",
         217 => x"03218100",
         218 => x"83204100",
         219 => x"13010108",
         220 => x"73002030",
         221 => x"e3eef6f6",
         222 => x"37370000",
         223 => x"93972700",
         224 => x"1307c7b5",
         225 => x"b387e700",
         226 => x"83a70700",
         227 => x"67800700",
         228 => x"eff05fda",
         229 => x"03258102",
         230 => x"6ff0dff5",
         231 => x"eff09fe0",
         232 => x"03258102",
         233 => x"6ff01ff5",
         234 => x"eff0dfe1",
         235 => x"03258102",
         236 => x"6ff05ff4",
         237 => x"eff01fe3",
         238 => x"03258102",
         239 => x"6ff09ff3",
         240 => x"eff01fdc",
         241 => x"03258102",
         242 => x"6ff0dff2",
         243 => x"9307600d",
         244 => x"6384f806",
         245 => x"9307900a",
         246 => x"6388f818",
         247 => x"63ca170f",
         248 => x"938878fc",
         249 => x"93074002",
         250 => x"63ec1703",
         251 => x"b7370000",
         252 => x"9387c7b8",
         253 => x"93982800",
         254 => x"b388f800",
         255 => x"83a70800",
         256 => x"67800700",
         257 => x"13050100",
         258 => x"eff01fc9",
         259 => x"03258102",
         260 => x"6ff05fee",
         261 => x"eff0dfce",
         262 => x"03258102",
         263 => x"6ff09fed",
         264 => x"ef104024",
         265 => x"93078005",
         266 => x"2320f500",
         267 => x"9307f0ff",
         268 => x"13850700",
         269 => x"6ff01fec",
         270 => x"63120510",
         271 => x"13858189",
         272 => x"13050500",
         273 => x"6ff01feb",
         274 => x"b7270000",
         275 => x"23a2f500",
         276 => x"93070000",
         277 => x"13850700",
         278 => x"6ff0dfe9",
         279 => x"93070000",
         280 => x"13850700",
         281 => x"6ff01fe9",
         282 => x"ef10c01f",
         283 => x"93079000",
         284 => x"2320f500",
         285 => x"9307f0ff",
         286 => x"13850700",
         287 => x"6ff09fe7",
         288 => x"13090600",
         289 => x"13840500",
         290 => x"635cc000",
         291 => x"b384c500",
         292 => x"03450400",
         293 => x"13041400",
         294 => x"eff05fbe",
         295 => x"e39a84fe",
         296 => x"13050900",
         297 => x"6ff01fe5",
         298 => x"13090600",
         299 => x"13840500",
         300 => x"e358c0fe",
         301 => x"b384c500",
         302 => x"eff01fbc",
         303 => x"2300a400",
         304 => x"13041400",
         305 => x"e31a94fe",
         306 => x"13050900",
         307 => x"6ff09fe2",
         308 => x"938808c0",
         309 => x"9307f000",
         310 => x"e3e417f5",
         311 => x"b7370000",
         312 => x"938707c2",
         313 => x"93982800",
         314 => x"b388f800",
         315 => x"83a70800",
         316 => x"67800700",
         317 => x"ef100017",
         318 => x"9307d000",
         319 => x"2320f500",
         320 => x"9307f0ff",
         321 => x"13850700",
         322 => x"6ff0dfde",
         323 => x"ef108015",
         324 => x"93072000",
         325 => x"2320f500",
         326 => x"9307f0ff",
         327 => x"13850700",
         328 => x"6ff05fdd",
         329 => x"ef100014",
         330 => x"9307f001",
         331 => x"2320f500",
         332 => x"9307f0ff",
         333 => x"13850700",
         334 => x"6ff0dfdb",
         335 => x"b7870020",
         336 => x"93870700",
         337 => x"13070040",
         338 => x"b387e740",
         339 => x"e36af5ee",
         340 => x"ef104011",
         341 => x"9307c000",
         342 => x"2320f500",
         343 => x"1305f0ff",
         344 => x"13050500",
         345 => x"6ff01fd9",
         346 => x"13090000",
         347 => x"93040500",
         348 => x"13040900",
         349 => x"93090900",
         350 => x"93070900",
         351 => x"732410c8",
         352 => x"f32910c0",
         353 => x"f32710c8",
         354 => x"e31af4fe",
         355 => x"37460f00",
         356 => x"13060624",
         357 => x"93060000",
         358 => x"13850900",
         359 => x"93050400",
         360 => x"ef005016",
         361 => x"37460f00",
         362 => x"23a4a400",
         363 => x"13060624",
         364 => x"93060000",
         365 => x"13850900",
         366 => x"93050400",
         367 => x"ef008051",
         368 => x"23a0a400",
         369 => x"23a2b400",
         370 => x"13050900",
         371 => x"6ff09fd2",
         372 => x"370700f0",
         373 => x"8327c702",
         374 => x"93f74700",
         375 => x"e38c07fe",
         376 => x"03250702",
         377 => x"1375f50f",
         378 => x"67800000",
         379 => x"b70700f0",
         380 => x"23a2a702",
         381 => x"23a4b702",
         382 => x"67800000",
         383 => x"1375f50f",
         384 => x"b70700f0",
         385 => x"23a0a702",
         386 => x"370700f0",
         387 => x"8327c702",
         388 => x"93f70701",
         389 => x"e38c07fe",
         390 => x"67800000",
         391 => x"630e0502",
         392 => x"130101ff",
         393 => x"23248100",
         394 => x"23261100",
         395 => x"13040500",
         396 => x"03450500",
         397 => x"630a0500",
         398 => x"13041400",
         399 => x"eff01ffc",
         400 => x"03450400",
         401 => x"e31a05fe",
         402 => x"8320c100",
         403 => x"03248100",
         404 => x"13010101",
         405 => x"67800000",
         406 => x"67800000",
         407 => x"13030500",
         408 => x"138e0500",
         409 => x"93080000",
         410 => x"63dc0500",
         411 => x"b337a000",
         412 => x"330eb040",
         413 => x"330efe40",
         414 => x"3303a040",
         415 => x"9308f0ff",
         416 => x"63dc0600",
         417 => x"b337c000",
         418 => x"b306d040",
         419 => x"93c8f8ff",
         420 => x"b386f640",
         421 => x"3306c040",
         422 => x"13070600",
         423 => x"13080300",
         424 => x"93070e00",
         425 => x"639c0628",
         426 => x"b7350000",
         427 => x"938505c6",
         428 => x"6376ce0e",
         429 => x"b7060100",
         430 => x"6378d60c",
         431 => x"93360610",
         432 => x"93c61600",
         433 => x"93963600",
         434 => x"3355d600",
         435 => x"b385a500",
         436 => x"83c50500",
         437 => x"13050002",
         438 => x"b386d500",
         439 => x"b305d540",
         440 => x"630cd500",
         441 => x"b317be00",
         442 => x"b356d300",
         443 => x"3317b600",
         444 => x"b3e7f600",
         445 => x"3318b300",
         446 => x"93550701",
         447 => x"33deb702",
         448 => x"13160701",
         449 => x"13560601",
         450 => x"b3f7b702",
         451 => x"13050e00",
         452 => x"3303c603",
         453 => x"93960701",
         454 => x"93570801",
         455 => x"b3e7d700",
         456 => x"63fe6700",
         457 => x"b307f700",
         458 => x"1305feff",
         459 => x"63e8e700",
         460 => x"63f66700",
         461 => x"1305eeff",
         462 => x"b387e700",
         463 => x"b3876740",
         464 => x"33d3b702",
         465 => x"13180801",
         466 => x"13580801",
         467 => x"b3f7b702",
         468 => x"b3066602",
         469 => x"93970701",
         470 => x"3368f800",
         471 => x"93070300",
         472 => x"637cd800",
         473 => x"33080701",
         474 => x"9307f3ff",
         475 => x"6366e800",
         476 => x"6374d800",
         477 => x"9307e3ff",
         478 => x"13150501",
         479 => x"3365f500",
         480 => x"93050000",
         481 => x"6f00000e",
         482 => x"37050001",
         483 => x"93060001",
         484 => x"e36ca6f2",
         485 => x"93068001",
         486 => x"6ff01ff3",
         487 => x"93060000",
         488 => x"630c0600",
         489 => x"b7070100",
         490 => x"637af60c",
         491 => x"93360610",
         492 => x"93c61600",
         493 => x"93963600",
         494 => x"b357d600",
         495 => x"b385f500",
         496 => x"83c70500",
         497 => x"b387d700",
         498 => x"93060002",
         499 => x"b385f640",
         500 => x"6390f60c",
         501 => x"b307ce40",
         502 => x"93051000",
         503 => x"13530701",
         504 => x"b3de6702",
         505 => x"13160701",
         506 => x"13560601",
         507 => x"93560801",
         508 => x"b3f76702",
         509 => x"13850e00",
         510 => x"330ed603",
         511 => x"93970701",
         512 => x"b3e7f600",
         513 => x"63fec701",
         514 => x"b307f700",
         515 => x"1385feff",
         516 => x"63e8e700",
         517 => x"63f6c701",
         518 => x"1385eeff",
         519 => x"b387e700",
         520 => x"b387c741",
         521 => x"33de6702",
         522 => x"13180801",
         523 => x"13580801",
         524 => x"b3f76702",
         525 => x"b306c603",
         526 => x"93970701",
         527 => x"3368f800",
         528 => x"93070e00",
         529 => x"637cd800",
         530 => x"33080701",
         531 => x"9307feff",
         532 => x"6366e800",
         533 => x"6374d800",
         534 => x"9307eeff",
         535 => x"13150501",
         536 => x"3365f500",
         537 => x"638a0800",
         538 => x"b337a000",
         539 => x"b305b040",
         540 => x"b385f540",
         541 => x"3305a040",
         542 => x"67800000",
         543 => x"b7070001",
         544 => x"93060001",
         545 => x"e36af6f2",
         546 => x"93068001",
         547 => x"6ff0dff2",
         548 => x"3317b600",
         549 => x"b356fe00",
         550 => x"13550701",
         551 => x"331ebe00",
         552 => x"b357f300",
         553 => x"b3e7c701",
         554 => x"33dea602",
         555 => x"13160701",
         556 => x"13560601",
         557 => x"3318b300",
         558 => x"b3f6a602",
         559 => x"3303c603",
         560 => x"93950601",
         561 => x"93d60701",
         562 => x"b3e6b600",
         563 => x"93050e00",
         564 => x"63fe6600",
         565 => x"b306d700",
         566 => x"9305feff",
         567 => x"63e8e600",
         568 => x"63f66600",
         569 => x"9305eeff",
         570 => x"b386e600",
         571 => x"b3866640",
         572 => x"33d3a602",
         573 => x"93970701",
         574 => x"93d70701",
         575 => x"b3f6a602",
         576 => x"33066602",
         577 => x"93960601",
         578 => x"b3e7d700",
         579 => x"93060300",
         580 => x"63fec700",
         581 => x"b307f700",
         582 => x"9306f3ff",
         583 => x"63e8e700",
         584 => x"63f6c700",
         585 => x"9306e3ff",
         586 => x"b387e700",
         587 => x"93950501",
         588 => x"b387c740",
         589 => x"b3e5d500",
         590 => x"6ff05fea",
         591 => x"6366de18",
         592 => x"b7070100",
         593 => x"63f4f604",
         594 => x"13b70610",
         595 => x"13471700",
         596 => x"13173700",
         597 => x"b7370000",
         598 => x"b3d5e600",
         599 => x"938707c6",
         600 => x"b387b700",
         601 => x"83c70700",
         602 => x"b387e700",
         603 => x"13070002",
         604 => x"b305f740",
         605 => x"6316f702",
         606 => x"13051000",
         607 => x"e3e4c6ef",
         608 => x"3335c300",
         609 => x"13451500",
         610 => x"6ff0dfed",
         611 => x"b7070001",
         612 => x"13070001",
         613 => x"e3e0f6fc",
         614 => x"13078001",
         615 => x"6ff09ffb",
         616 => x"3357f600",
         617 => x"b396b600",
         618 => x"b366d700",
         619 => x"3357fe00",
         620 => x"331ebe00",
         621 => x"b357f300",
         622 => x"b3e7c701",
         623 => x"13de0601",
         624 => x"335fc703",
         625 => x"13980601",
         626 => x"13580801",
         627 => x"3316b600",
         628 => x"3377c703",
         629 => x"b30ee803",
         630 => x"13150701",
         631 => x"13d70701",
         632 => x"3367a700",
         633 => x"13050f00",
         634 => x"637ed701",
         635 => x"3387e600",
         636 => x"1305ffff",
         637 => x"6368d700",
         638 => x"6376d701",
         639 => x"1305efff",
         640 => x"3307d700",
         641 => x"3307d741",
         642 => x"b35ec703",
         643 => x"93970701",
         644 => x"93d70701",
         645 => x"3377c703",
         646 => x"3308d803",
         647 => x"13170701",
         648 => x"b3e7e700",
         649 => x"13870e00",
         650 => x"63fe0701",
         651 => x"b387f600",
         652 => x"1387feff",
         653 => x"63e8d700",
         654 => x"63f60701",
         655 => x"1387eeff",
         656 => x"b387d700",
         657 => x"13150501",
         658 => x"b70e0100",
         659 => x"3365e500",
         660 => x"9386feff",
         661 => x"3377d500",
         662 => x"b3870741",
         663 => x"b376d600",
         664 => x"13580501",
         665 => x"13560601",
         666 => x"330ed702",
         667 => x"b306d802",
         668 => x"3307c702",
         669 => x"3308c802",
         670 => x"3306d700",
         671 => x"13570e01",
         672 => x"3307c700",
         673 => x"6374d700",
         674 => x"3308d801",
         675 => x"93560701",
         676 => x"b3860601",
         677 => x"63e6d702",
         678 => x"e394d7ce",
         679 => x"b7070100",
         680 => x"9387f7ff",
         681 => x"3377f700",
         682 => x"13170701",
         683 => x"337efe00",
         684 => x"3313b300",
         685 => x"3307c701",
         686 => x"93050000",
         687 => x"e374e3da",
         688 => x"1305f5ff",
         689 => x"6ff0dfcb",
         690 => x"93050000",
         691 => x"13050000",
         692 => x"6ff05fd9",
         693 => x"93080500",
         694 => x"13830500",
         695 => x"13070600",
         696 => x"13080500",
         697 => x"93870500",
         698 => x"63920628",
         699 => x"b7350000",
         700 => x"938505c6",
         701 => x"6376c30e",
         702 => x"b7060100",
         703 => x"6378d60c",
         704 => x"93360610",
         705 => x"93c61600",
         706 => x"93963600",
         707 => x"3355d600",
         708 => x"b385a500",
         709 => x"83c50500",
         710 => x"13050002",
         711 => x"b386d500",
         712 => x"b305d540",
         713 => x"630cd500",
         714 => x"b317b300",
         715 => x"b3d6d800",
         716 => x"3317b600",
         717 => x"b3e7f600",
         718 => x"3398b800",
         719 => x"93550701",
         720 => x"33d3b702",
         721 => x"13160701",
         722 => x"13560601",
         723 => x"b3f7b702",
         724 => x"13050300",
         725 => x"b3086602",
         726 => x"93960701",
         727 => x"93570801",
         728 => x"b3e7d700",
         729 => x"63fe1701",
         730 => x"b307f700",
         731 => x"1305f3ff",
         732 => x"63e8e700",
         733 => x"63f61701",
         734 => x"1305e3ff",
         735 => x"b387e700",
         736 => x"b3871741",
         737 => x"b3d8b702",
         738 => x"13180801",
         739 => x"13580801",
         740 => x"b3f7b702",
         741 => x"b3061603",
         742 => x"93970701",
         743 => x"3368f800",
         744 => x"93870800",
         745 => x"637cd800",
         746 => x"33080701",
         747 => x"9387f8ff",
         748 => x"6366e800",
         749 => x"6374d800",
         750 => x"9387e8ff",
         751 => x"13150501",
         752 => x"3365f500",
         753 => x"93050000",
         754 => x"67800000",
         755 => x"37050001",
         756 => x"93060001",
         757 => x"e36ca6f2",
         758 => x"93068001",
         759 => x"6ff01ff3",
         760 => x"93060000",
         761 => x"630c0600",
         762 => x"b7070100",
         763 => x"6370f60c",
         764 => x"93360610",
         765 => x"93c61600",
         766 => x"93963600",
         767 => x"b357d600",
         768 => x"b385f500",
         769 => x"83c70500",
         770 => x"b387d700",
         771 => x"93060002",
         772 => x"b385f640",
         773 => x"6396f60a",
         774 => x"b307c340",
         775 => x"93051000",
         776 => x"93580701",
         777 => x"33de1703",
         778 => x"13160701",
         779 => x"13560601",
         780 => x"93560801",
         781 => x"b3f71703",
         782 => x"13050e00",
         783 => x"3303c603",
         784 => x"93970701",
         785 => x"b3e7f600",
         786 => x"63fe6700",
         787 => x"b307f700",
         788 => x"1305feff",
         789 => x"63e8e700",
         790 => x"63f66700",
         791 => x"1305eeff",
         792 => x"b387e700",
         793 => x"b3876740",
         794 => x"33d31703",
         795 => x"13180801",
         796 => x"13580801",
         797 => x"b3f71703",
         798 => x"b3066602",
         799 => x"93970701",
         800 => x"3368f800",
         801 => x"93070300",
         802 => x"637cd800",
         803 => x"33080701",
         804 => x"9307f3ff",
         805 => x"6366e800",
         806 => x"6374d800",
         807 => x"9307e3ff",
         808 => x"13150501",
         809 => x"3365f500",
         810 => x"67800000",
         811 => x"b7070001",
         812 => x"93060001",
         813 => x"e364f6f4",
         814 => x"93068001",
         815 => x"6ff01ff4",
         816 => x"3317b600",
         817 => x"b356f300",
         818 => x"13550701",
         819 => x"3313b300",
         820 => x"b3d7f800",
         821 => x"b3e76700",
         822 => x"33d3a602",
         823 => x"13160701",
         824 => x"13560601",
         825 => x"3398b800",
         826 => x"b3f6a602",
         827 => x"b3086602",
         828 => x"93950601",
         829 => x"93d60701",
         830 => x"b3e6b600",
         831 => x"93050300",
         832 => x"63fe1601",
         833 => x"b306d700",
         834 => x"9305f3ff",
         835 => x"63e8e600",
         836 => x"63f61601",
         837 => x"9305e3ff",
         838 => x"b386e600",
         839 => x"b3861641",
         840 => x"b3d8a602",
         841 => x"93970701",
         842 => x"93d70701",
         843 => x"b3f6a602",
         844 => x"33061603",
         845 => x"93960601",
         846 => x"b3e7d700",
         847 => x"93860800",
         848 => x"63fec700",
         849 => x"b307f700",
         850 => x"9386f8ff",
         851 => x"63e8e700",
         852 => x"63f6c700",
         853 => x"9386e8ff",
         854 => x"b387e700",
         855 => x"93950501",
         856 => x"b387c740",
         857 => x"b3e5d500",
         858 => x"6ff09feb",
         859 => x"63e6d518",
         860 => x"b7070100",
         861 => x"63f4f604",
         862 => x"13b70610",
         863 => x"13471700",
         864 => x"13173700",
         865 => x"b7370000",
         866 => x"b3d5e600",
         867 => x"938707c6",
         868 => x"b387b700",
         869 => x"83c70700",
         870 => x"b387e700",
         871 => x"13070002",
         872 => x"b305f740",
         873 => x"6316f702",
         874 => x"13051000",
         875 => x"e3ee66e0",
         876 => x"33b5c800",
         877 => x"13451500",
         878 => x"67800000",
         879 => x"b7070001",
         880 => x"13070001",
         881 => x"e3e0f6fc",
         882 => x"13078001",
         883 => x"6ff09ffb",
         884 => x"3357f600",
         885 => x"b396b600",
         886 => x"b366d700",
         887 => x"3357f300",
         888 => x"3313b300",
         889 => x"b3d7f800",
         890 => x"b3e76700",
         891 => x"13d30601",
         892 => x"b35e6702",
         893 => x"13980601",
         894 => x"13580801",
         895 => x"3316b600",
         896 => x"33776702",
         897 => x"330ed803",
         898 => x"13150701",
         899 => x"13d70701",
         900 => x"3367a700",
         901 => x"13850e00",
         902 => x"637ec701",
         903 => x"3387e600",
         904 => x"1385feff",
         905 => x"6368d700",
         906 => x"6376c701",
         907 => x"1385eeff",
         908 => x"3307d700",
         909 => x"3307c741",
         910 => x"335e6702",
         911 => x"93970701",
         912 => x"93d70701",
         913 => x"33776702",
         914 => x"3308c803",
         915 => x"13170701",
         916 => x"b3e7e700",
         917 => x"13070e00",
         918 => x"63fe0701",
         919 => x"b387f600",
         920 => x"1307feff",
         921 => x"63e8d700",
         922 => x"63f60701",
         923 => x"1307eeff",
         924 => x"b387d700",
         925 => x"13150501",
         926 => x"370e0100",
         927 => x"3365e500",
         928 => x"9306feff",
         929 => x"3377d500",
         930 => x"b3870741",
         931 => x"b376d600",
         932 => x"13580501",
         933 => x"13560601",
         934 => x"3303d702",
         935 => x"b306d802",
         936 => x"3307c702",
         937 => x"3308c802",
         938 => x"3306d700",
         939 => x"13570301",
         940 => x"3307c700",
         941 => x"6374d700",
         942 => x"3308c801",
         943 => x"93560701",
         944 => x"b3860601",
         945 => x"63e6d702",
         946 => x"e39ed7ce",
         947 => x"b7070100",
         948 => x"9387f7ff",
         949 => x"3377f700",
         950 => x"13170701",
         951 => x"3373f300",
         952 => x"b398b800",
         953 => x"33076700",
         954 => x"93050000",
         955 => x"e3fee8cc",
         956 => x"1305f5ff",
         957 => x"6ff01fcd",
         958 => x"93050000",
         959 => x"13050000",
         960 => x"67800000",
         961 => x"13080600",
         962 => x"93070500",
         963 => x"13870500",
         964 => x"63960620",
         965 => x"b7380000",
         966 => x"938808c6",
         967 => x"63fcc50c",
         968 => x"b7060100",
         969 => x"637ed60a",
         970 => x"93360610",
         971 => x"93c61600",
         972 => x"93963600",
         973 => x"3353d600",
         974 => x"b3886800",
         975 => x"83c80800",
         976 => x"13030002",
         977 => x"b386d800",
         978 => x"b308d340",
         979 => x"630cd300",
         980 => x"33971501",
         981 => x"b356d500",
         982 => x"33181601",
         983 => x"33e7e600",
         984 => x"b3171501",
         985 => x"13560801",
         986 => x"b356c702",
         987 => x"13150801",
         988 => x"13550501",
         989 => x"3377c702",
         990 => x"b386a602",
         991 => x"93150701",
         992 => x"13d70701",
         993 => x"3367b700",
         994 => x"637ad700",
         995 => x"3307e800",
         996 => x"63660701",
         997 => x"6374d700",
         998 => x"33070701",
         999 => x"3307d740",
        1000 => x"b356c702",
        1001 => x"3377c702",
        1002 => x"b386a602",
        1003 => x"93970701",
        1004 => x"13170701",
        1005 => x"93d70701",
        1006 => x"b3e7e700",
        1007 => x"63fad700",
        1008 => x"b307f800",
        1009 => x"63e60701",
        1010 => x"63f4d700",
        1011 => x"b3870701",
        1012 => x"b387d740",
        1013 => x"33d51701",
        1014 => x"93050000",
        1015 => x"67800000",
        1016 => x"37030001",
        1017 => x"93060001",
        1018 => x"e36666f4",
        1019 => x"93068001",
        1020 => x"6ff05ff4",
        1021 => x"93060000",
        1022 => x"630c0600",
        1023 => x"37070100",
        1024 => x"637ee606",
        1025 => x"93360610",
        1026 => x"93c61600",
        1027 => x"93963600",
        1028 => x"3357d600",
        1029 => x"b388e800",
        1030 => x"03c70800",
        1031 => x"3307d700",
        1032 => x"93060002",
        1033 => x"b388e640",
        1034 => x"6394e606",
        1035 => x"3387c540",
        1036 => x"93550801",
        1037 => x"3356b702",
        1038 => x"13150801",
        1039 => x"13550501",
        1040 => x"93d60701",
        1041 => x"3377b702",
        1042 => x"3306a602",
        1043 => x"13170701",
        1044 => x"33e7e600",
        1045 => x"637ac700",
        1046 => x"3307e800",
        1047 => x"63660701",
        1048 => x"6374c700",
        1049 => x"33070701",
        1050 => x"3307c740",
        1051 => x"b356b702",
        1052 => x"3377b702",
        1053 => x"b386a602",
        1054 => x"6ff05ff3",
        1055 => x"37070001",
        1056 => x"93060001",
        1057 => x"e366e6f8",
        1058 => x"93068001",
        1059 => x"6ff05ff8",
        1060 => x"33181601",
        1061 => x"b3d6e500",
        1062 => x"b3171501",
        1063 => x"b3951501",
        1064 => x"3357e500",
        1065 => x"13550801",
        1066 => x"3367b700",
        1067 => x"b3d5a602",
        1068 => x"13130801",
        1069 => x"13530301",
        1070 => x"b3f6a602",
        1071 => x"b3856502",
        1072 => x"13960601",
        1073 => x"93560701",
        1074 => x"b3e6c600",
        1075 => x"63fab600",
        1076 => x"b306d800",
        1077 => x"63e60601",
        1078 => x"63f4b600",
        1079 => x"b3860601",
        1080 => x"b386b640",
        1081 => x"33d6a602",
        1082 => x"13170701",
        1083 => x"13570701",
        1084 => x"b3f6a602",
        1085 => x"33066602",
        1086 => x"93960601",
        1087 => x"3367d700",
        1088 => x"637ac700",
        1089 => x"3307e800",
        1090 => x"63660701",
        1091 => x"6374c700",
        1092 => x"33070701",
        1093 => x"3307c740",
        1094 => x"6ff09ff1",
        1095 => x"63e4d51c",
        1096 => x"37080100",
        1097 => x"63fe0605",
        1098 => x"13b80610",
        1099 => x"13481800",
        1100 => x"13183800",
        1101 => x"b7380000",
        1102 => x"33d30601",
        1103 => x"938808c6",
        1104 => x"b3886800",
        1105 => x"83c80800",
        1106 => x"13030002",
        1107 => x"b3880801",
        1108 => x"33081341",
        1109 => x"63101305",
        1110 => x"63e4b600",
        1111 => x"636cc500",
        1112 => x"3306c540",
        1113 => x"b386d540",
        1114 => x"3337c500",
        1115 => x"93070600",
        1116 => x"3387e640",
        1117 => x"13850700",
        1118 => x"93050700",
        1119 => x"67800000",
        1120 => x"b7080001",
        1121 => x"13080001",
        1122 => x"e3e616fb",
        1123 => x"13088001",
        1124 => x"6ff05ffa",
        1125 => x"b3571601",
        1126 => x"b3960601",
        1127 => x"b3e6d700",
        1128 => x"33d71501",
        1129 => x"13de0601",
        1130 => x"335fc703",
        1131 => x"13930601",
        1132 => x"13530301",
        1133 => x"b3970501",
        1134 => x"b3551501",
        1135 => x"b3e5f500",
        1136 => x"93d70501",
        1137 => x"33160601",
        1138 => x"33150501",
        1139 => x"3377c703",
        1140 => x"b30ee303",
        1141 => x"13170701",
        1142 => x"b3e7e700",
        1143 => x"13070f00",
        1144 => x"63fed701",
        1145 => x"b387f600",
        1146 => x"1307ffff",
        1147 => x"63e8d700",
        1148 => x"63f6d701",
        1149 => x"1307efff",
        1150 => x"b387d700",
        1151 => x"b387d741",
        1152 => x"b3dec703",
        1153 => x"93950501",
        1154 => x"93d50501",
        1155 => x"b3f7c703",
        1156 => x"138e0e00",
        1157 => x"3303d303",
        1158 => x"93970701",
        1159 => x"b3e5f500",
        1160 => x"63fe6500",
        1161 => x"b385b600",
        1162 => x"138efeff",
        1163 => x"63e8d500",
        1164 => x"63f66500",
        1165 => x"138eeeff",
        1166 => x"b385d500",
        1167 => x"93170701",
        1168 => x"370f0100",
        1169 => x"b3e7c701",
        1170 => x"b3856540",
        1171 => x"1303ffff",
        1172 => x"33f76700",
        1173 => x"135e0601",
        1174 => x"93d70701",
        1175 => x"33736600",
        1176 => x"b30e6702",
        1177 => x"33836702",
        1178 => x"3307c703",
        1179 => x"b387c703",
        1180 => x"330e6700",
        1181 => x"13d70e01",
        1182 => x"3307c701",
        1183 => x"63746700",
        1184 => x"b387e701",
        1185 => x"13530701",
        1186 => x"b307f300",
        1187 => x"37030100",
        1188 => x"1303f3ff",
        1189 => x"33776700",
        1190 => x"13170701",
        1191 => x"b3fe6e00",
        1192 => x"3307d701",
        1193 => x"63e6f500",
        1194 => x"639ef500",
        1195 => x"637ce500",
        1196 => x"3306c740",
        1197 => x"3333c700",
        1198 => x"b306d300",
        1199 => x"13070600",
        1200 => x"b387d740",
        1201 => x"3307e540",
        1202 => x"3335e500",
        1203 => x"b385f540",
        1204 => x"b385a540",
        1205 => x"b3981501",
        1206 => x"33570701",
        1207 => x"33e5e800",
        1208 => x"b3d50501",
        1209 => x"67800000",
        1210 => x"13030500",
        1211 => x"630e0600",
        1212 => x"83830500",
        1213 => x"23007300",
        1214 => x"1306f6ff",
        1215 => x"13031300",
        1216 => x"93851500",
        1217 => x"e31606fe",
        1218 => x"67800000",
        1219 => x"13030500",
        1220 => x"630a0600",
        1221 => x"2300b300",
        1222 => x"1306f6ff",
        1223 => x"13031300",
        1224 => x"e31a06fe",
        1225 => x"67800000",
        1226 => x"630c0602",
        1227 => x"13030500",
        1228 => x"93061000",
        1229 => x"636ab500",
        1230 => x"9306f0ff",
        1231 => x"1307f6ff",
        1232 => x"3303e300",
        1233 => x"b385e500",
        1234 => x"83830500",
        1235 => x"23007300",
        1236 => x"1306f6ff",
        1237 => x"3303d300",
        1238 => x"b385d500",
        1239 => x"e31606fe",
        1240 => x"67800000",
        1241 => x"130101f9",
        1242 => x"23248106",
        1243 => x"23229106",
        1244 => x"23261106",
        1245 => x"23202107",
        1246 => x"232e3105",
        1247 => x"232c4105",
        1248 => x"232a5105",
        1249 => x"23286105",
        1250 => x"23267105",
        1251 => x"23248105",
        1252 => x"23229105",
        1253 => x"2320a105",
        1254 => x"93040500",
        1255 => x"13840500",
        1256 => x"232c0100",
        1257 => x"232e0100",
        1258 => x"23200102",
        1259 => x"23220102",
        1260 => x"23240102",
        1261 => x"23260102",
        1262 => x"23280102",
        1263 => x"232a0102",
        1264 => x"232c0102",
        1265 => x"232e0102",
        1266 => x"97f2ffff",
        1267 => x"938202e5",
        1268 => x"73905230",
        1269 => x"93050004",
        1270 => x"1305101b",
        1271 => x"eff00fa1",
        1272 => x"37877d01",
        1273 => x"b70700f0",
        1274 => x"1307f783",
        1275 => x"23a6e708",
        1276 => x"93061001",
        1277 => x"37170000",
        1278 => x"23a0d708",
        1279 => x"13077738",
        1280 => x"23a8e70a",
        1281 => x"37270000",
        1282 => x"1307f770",
        1283 => x"23a6e70a",
        1284 => x"23a0d70a",
        1285 => x"13078070",
        1286 => x"23a0e706",
        1287 => x"3707f900",
        1288 => x"13078700",
        1289 => x"23a0e704",
        1290 => x"93020008",
        1291 => x"73904230",
        1292 => x"b7220000",
        1293 => x"93828280",
        1294 => x"73900230",
        1295 => x"b7390000",
        1296 => x"138509da",
        1297 => x"eff08f9d",
        1298 => x"63549002",
        1299 => x"1389f4ff",
        1300 => x"9304f0ff",
        1301 => x"03250400",
        1302 => x"1309f9ff",
        1303 => x"13044400",
        1304 => x"eff0cf9b",
        1305 => x"138509da",
        1306 => x"eff04f9b",
        1307 => x"e31499fe",
        1308 => x"37350000",
        1309 => x"b7faeeee",
        1310 => x"130545d7",
        1311 => x"b7090010",
        1312 => x"37140000",
        1313 => x"1389faee",
        1314 => x"eff04f99",
        1315 => x"373b0000",
        1316 => x"9389f9ff",
        1317 => x"938aeaee",
        1318 => x"130404e1",
        1319 => x"93040000",
        1320 => x"b71b0000",
        1321 => x"938b0b2c",
        1322 => x"130af000",
        1323 => x"93050000",
        1324 => x"13058100",
        1325 => x"ef008036",
        1326 => x"938bfbff",
        1327 => x"630a0502",
        1328 => x"e3960bfe",
        1329 => x"73001000",
        1330 => x"b70700f0",
        1331 => x"9306f00f",
        1332 => x"23a4d706",
        1333 => x"03a70704",
        1334 => x"93860704",
        1335 => x"13670730",
        1336 => x"23a0e704",
        1337 => x"93070009",
        1338 => x"23a4f600",
        1339 => x"6ff05ffb",
        1340 => x"032c8100",
        1341 => x"8325c100",
        1342 => x"13060400",
        1343 => x"9357cc01",
        1344 => x"13974500",
        1345 => x"b367f700",
        1346 => x"b3f73701",
        1347 => x"33773c01",
        1348 => x"13d5f541",
        1349 => x"13d88501",
        1350 => x"3307f700",
        1351 => x"33070701",
        1352 => x"9377d500",
        1353 => x"3307f700",
        1354 => x"33774703",
        1355 => x"937725ff",
        1356 => x"93860400",
        1357 => x"13050c00",
        1358 => x"3307f700",
        1359 => x"b307ec40",
        1360 => x"1357f741",
        1361 => x"3338fc00",
        1362 => x"3387e540",
        1363 => x"33070741",
        1364 => x"b3885703",
        1365 => x"33072703",
        1366 => x"33b82703",
        1367 => x"33071701",
        1368 => x"b3872703",
        1369 => x"33070701",
        1370 => x"1358f741",
        1371 => x"13783800",
        1372 => x"b307f800",
        1373 => x"33b80701",
        1374 => x"3307e800",
        1375 => x"1318e701",
        1376 => x"93d72700",
        1377 => x"b367f800",
        1378 => x"13582740",
        1379 => x"93184800",
        1380 => x"13d3c701",
        1381 => x"33e36800",
        1382 => x"33733301",
        1383 => x"b3f83701",
        1384 => x"135e8801",
        1385 => x"1357f741",
        1386 => x"b3886800",
        1387 => x"b388c801",
        1388 => x"1373d700",
        1389 => x"b3886800",
        1390 => x"b3f84803",
        1391 => x"137727ff",
        1392 => x"939c4700",
        1393 => x"b38cfc40",
        1394 => x"939c2c00",
        1395 => x"b30c9c41",
        1396 => x"b388e800",
        1397 => x"33871741",
        1398 => x"93d8f841",
        1399 => x"33b3e700",
        1400 => x"33081841",
        1401 => x"33086840",
        1402 => x"33082803",
        1403 => x"33035703",
        1404 => x"b3382703",
        1405 => x"33086800",
        1406 => x"33072703",
        1407 => x"33081801",
        1408 => x"9358f841",
        1409 => x"93f83800",
        1410 => x"3387e800",
        1411 => x"b3381701",
        1412 => x"b3880801",
        1413 => x"9398e801",
        1414 => x"13572700",
        1415 => x"33e7e800",
        1416 => x"13184700",
        1417 => x"3307e840",
        1418 => x"13172700",
        1419 => x"338de740",
        1420 => x"eff0cf82",
        1421 => x"83260101",
        1422 => x"13070500",
        1423 => x"13880c00",
        1424 => x"93070d00",
        1425 => x"13060c00",
        1426 => x"93054bda",
        1427 => x"13058101",
        1428 => x"ef00c015",
        1429 => x"13058101",
        1430 => x"efe05ffc",
        1431 => x"e3980be4",
        1432 => x"6ff05fe6",
        1433 => x"03a5c187",
        1434 => x"67800000",
        1435 => x"130101ff",
        1436 => x"23248100",
        1437 => x"23261100",
        1438 => x"93070000",
        1439 => x"13040500",
        1440 => x"63880700",
        1441 => x"93050000",
        1442 => x"97000000",
        1443 => x"e7000000",
        1444 => x"b7370000",
        1445 => x"03a547f0",
        1446 => x"83278502",
        1447 => x"63840700",
        1448 => x"e7800700",
        1449 => x"13050400",
        1450 => x"ef100035",
        1451 => x"130101ff",
        1452 => x"23248100",
        1453 => x"23229100",
        1454 => x"37340000",
        1455 => x"b7340000",
        1456 => x"938784f0",
        1457 => x"130484f0",
        1458 => x"3304f440",
        1459 => x"23202101",
        1460 => x"23261100",
        1461 => x"13542440",
        1462 => x"938484f0",
        1463 => x"13090000",
        1464 => x"63108904",
        1465 => x"b7340000",
        1466 => x"37340000",
        1467 => x"938784f0",
        1468 => x"130484f0",
        1469 => x"3304f440",
        1470 => x"13542440",
        1471 => x"938484f0",
        1472 => x"13090000",
        1473 => x"63188902",
        1474 => x"8320c100",
        1475 => x"03248100",
        1476 => x"83244100",
        1477 => x"03290100",
        1478 => x"13010101",
        1479 => x"67800000",
        1480 => x"83a70400",
        1481 => x"13091900",
        1482 => x"93844400",
        1483 => x"e7800700",
        1484 => x"6ff01ffb",
        1485 => x"83a70400",
        1486 => x"13091900",
        1487 => x"93844400",
        1488 => x"e7800700",
        1489 => x"6ff01ffc",
        1490 => x"130101f6",
        1491 => x"232af108",
        1492 => x"b7070080",
        1493 => x"93c7f7ff",
        1494 => x"232ef100",
        1495 => x"2328f100",
        1496 => x"b707ffff",
        1497 => x"2326d108",
        1498 => x"2324b100",
        1499 => x"232cb100",
        1500 => x"93878720",
        1501 => x"9306c108",
        1502 => x"93058100",
        1503 => x"232e1106",
        1504 => x"232af100",
        1505 => x"2328e108",
        1506 => x"232c0109",
        1507 => x"232e1109",
        1508 => x"2322d100",
        1509 => x"ef00c040",
        1510 => x"83278100",
        1511 => x"23800700",
        1512 => x"8320c107",
        1513 => x"1301010a",
        1514 => x"67800000",
        1515 => x"130101f6",
        1516 => x"232af108",
        1517 => x"b7070080",
        1518 => x"93c7f7ff",
        1519 => x"232ef100",
        1520 => x"2328f100",
        1521 => x"b707ffff",
        1522 => x"93878720",
        1523 => x"232af100",
        1524 => x"2324a100",
        1525 => x"232ca100",
        1526 => x"03a5c187",
        1527 => x"2324c108",
        1528 => x"2326d108",
        1529 => x"13860500",
        1530 => x"93068108",
        1531 => x"93058100",
        1532 => x"232e1106",
        1533 => x"2328e108",
        1534 => x"232c0109",
        1535 => x"232e1109",
        1536 => x"2322d100",
        1537 => x"ef00c039",
        1538 => x"83278100",
        1539 => x"23800700",
        1540 => x"8320c107",
        1541 => x"1301010a",
        1542 => x"67800000",
        1543 => x"13860500",
        1544 => x"93050500",
        1545 => x"03a5c187",
        1546 => x"6f004000",
        1547 => x"130101ff",
        1548 => x"23248100",
        1549 => x"23229100",
        1550 => x"13040500",
        1551 => x"13850500",
        1552 => x"93050600",
        1553 => x"23261100",
        1554 => x"23a20188",
        1555 => x"ef10c01d",
        1556 => x"9307f0ff",
        1557 => x"6318f500",
        1558 => x"83a74188",
        1559 => x"63840700",
        1560 => x"2320f400",
        1561 => x"8320c100",
        1562 => x"03248100",
        1563 => x"83244100",
        1564 => x"13010101",
        1565 => x"67800000",
        1566 => x"130101fe",
        1567 => x"23282101",
        1568 => x"03a98500",
        1569 => x"232c8100",
        1570 => x"23263101",
        1571 => x"23225101",
        1572 => x"23206101",
        1573 => x"232e1100",
        1574 => x"232a9100",
        1575 => x"23244101",
        1576 => x"83aa0500",
        1577 => x"13840500",
        1578 => x"130b0600",
        1579 => x"93890600",
        1580 => x"63ec2609",
        1581 => x"8397c500",
        1582 => x"13f70748",
        1583 => x"63040708",
        1584 => x"03274401",
        1585 => x"93043000",
        1586 => x"83a50501",
        1587 => x"b384e402",
        1588 => x"13072000",
        1589 => x"b38aba40",
        1590 => x"130a0500",
        1591 => x"b3c4e402",
        1592 => x"13871600",
        1593 => x"33075701",
        1594 => x"63f4e400",
        1595 => x"93040700",
        1596 => x"93f70740",
        1597 => x"6386070a",
        1598 => x"93850400",
        1599 => x"13050a00",
        1600 => x"ef001067",
        1601 => x"13090500",
        1602 => x"630c050a",
        1603 => x"83250401",
        1604 => x"13860a00",
        1605 => x"eff05f9d",
        1606 => x"8357c400",
        1607 => x"93f7f7b7",
        1608 => x"93e70708",
        1609 => x"2316f400",
        1610 => x"23282401",
        1611 => x"232a9400",
        1612 => x"33095901",
        1613 => x"b3845441",
        1614 => x"23202401",
        1615 => x"23249400",
        1616 => x"13890900",
        1617 => x"63f42901",
        1618 => x"13890900",
        1619 => x"03250400",
        1620 => x"13060900",
        1621 => x"93050b00",
        1622 => x"eff01f9d",
        1623 => x"83278400",
        1624 => x"13050000",
        1625 => x"b3872741",
        1626 => x"2324f400",
        1627 => x"83270400",
        1628 => x"b3872701",
        1629 => x"2320f400",
        1630 => x"8320c101",
        1631 => x"03248101",
        1632 => x"83244101",
        1633 => x"03290101",
        1634 => x"8329c100",
        1635 => x"032a8100",
        1636 => x"832a4100",
        1637 => x"032b0100",
        1638 => x"13010102",
        1639 => x"67800000",
        1640 => x"13860400",
        1641 => x"13050a00",
        1642 => x"ef001071",
        1643 => x"13090500",
        1644 => x"e31c05f6",
        1645 => x"83250401",
        1646 => x"13050a00",
        1647 => x"ef00d04b",
        1648 => x"9307c000",
        1649 => x"2320fa00",
        1650 => x"8357c400",
        1651 => x"1305f0ff",
        1652 => x"93e70704",
        1653 => x"2316f400",
        1654 => x"6ff01ffa",
        1655 => x"83278600",
        1656 => x"130101fd",
        1657 => x"232e3101",
        1658 => x"23286101",
        1659 => x"23261102",
        1660 => x"23248102",
        1661 => x"23229102",
        1662 => x"23202103",
        1663 => x"232c4101",
        1664 => x"232a5101",
        1665 => x"23267101",
        1666 => x"23248101",
        1667 => x"23229101",
        1668 => x"2320a101",
        1669 => x"032b0600",
        1670 => x"93090600",
        1671 => x"63940712",
        1672 => x"13050000",
        1673 => x"8320c102",
        1674 => x"03248102",
        1675 => x"23a20900",
        1676 => x"83244102",
        1677 => x"03290102",
        1678 => x"8329c101",
        1679 => x"032a8101",
        1680 => x"832a4101",
        1681 => x"032b0101",
        1682 => x"832bc100",
        1683 => x"032c8100",
        1684 => x"832c4100",
        1685 => x"032d0100",
        1686 => x"13010103",
        1687 => x"67800000",
        1688 => x"832b0b00",
        1689 => x"032d4b00",
        1690 => x"130b8b00",
        1691 => x"03298400",
        1692 => x"832a0400",
        1693 => x"e3060dfe",
        1694 => x"63642d09",
        1695 => x"8317c400",
        1696 => x"13f70748",
        1697 => x"630e0706",
        1698 => x"83244401",
        1699 => x"83250401",
        1700 => x"b3049c02",
        1701 => x"b38aba40",
        1702 => x"13871a00",
        1703 => x"3307a701",
        1704 => x"b3c49403",
        1705 => x"63f4e400",
        1706 => x"93040700",
        1707 => x"93f70740",
        1708 => x"6388070a",
        1709 => x"93850400",
        1710 => x"13050a00",
        1711 => x"ef00504b",
        1712 => x"13090500",
        1713 => x"630e050a",
        1714 => x"83250401",
        1715 => x"13860a00",
        1716 => x"eff09f81",
        1717 => x"8357c400",
        1718 => x"93f7f7b7",
        1719 => x"93e70708",
        1720 => x"2316f400",
        1721 => x"23282401",
        1722 => x"232a9400",
        1723 => x"33095901",
        1724 => x"b3845441",
        1725 => x"23202401",
        1726 => x"23249400",
        1727 => x"13090d00",
        1728 => x"63742d01",
        1729 => x"13090d00",
        1730 => x"03250400",
        1731 => x"13060900",
        1732 => x"93850b00",
        1733 => x"eff05f81",
        1734 => x"83278400",
        1735 => x"b3872741",
        1736 => x"2324f400",
        1737 => x"83270400",
        1738 => x"b3872701",
        1739 => x"2320f400",
        1740 => x"83a78900",
        1741 => x"b387a741",
        1742 => x"23a4f900",
        1743 => x"e39207f2",
        1744 => x"6ff01fee",
        1745 => x"130a0500",
        1746 => x"13840500",
        1747 => x"930b0000",
        1748 => x"130d0000",
        1749 => x"130c3000",
        1750 => x"930c2000",
        1751 => x"6ff01ff1",
        1752 => x"13860400",
        1753 => x"13050a00",
        1754 => x"ef001055",
        1755 => x"13090500",
        1756 => x"e31a05f6",
        1757 => x"83250401",
        1758 => x"13050a00",
        1759 => x"ef00d02f",
        1760 => x"9307c000",
        1761 => x"2320fa00",
        1762 => x"8357c400",
        1763 => x"1305f0ff",
        1764 => x"93e70704",
        1765 => x"2316f400",
        1766 => x"23a40900",
        1767 => x"6ff09fe8",
        1768 => x"83d7c500",
        1769 => x"130101f5",
        1770 => x"2324810a",
        1771 => x"2322910a",
        1772 => x"2320210b",
        1773 => x"232c4109",
        1774 => x"2326110a",
        1775 => x"232e3109",
        1776 => x"232a5109",
        1777 => x"23286109",
        1778 => x"23267109",
        1779 => x"23248109",
        1780 => x"23229109",
        1781 => x"2320a109",
        1782 => x"232eb107",
        1783 => x"93f70708",
        1784 => x"130a0500",
        1785 => x"13890500",
        1786 => x"93040600",
        1787 => x"13840600",
        1788 => x"63880706",
        1789 => x"83a70501",
        1790 => x"63940706",
        1791 => x"93050004",
        1792 => x"ef001037",
        1793 => x"2320a900",
        1794 => x"2328a900",
        1795 => x"63160504",
        1796 => x"9307c000",
        1797 => x"2320fa00",
        1798 => x"1305f0ff",
        1799 => x"8320c10a",
        1800 => x"0324810a",
        1801 => x"8324410a",
        1802 => x"0329010a",
        1803 => x"8329c109",
        1804 => x"032a8109",
        1805 => x"832a4109",
        1806 => x"032b0109",
        1807 => x"832bc108",
        1808 => x"032c8108",
        1809 => x"832c4108",
        1810 => x"032d0108",
        1811 => x"832dc107",
        1812 => x"1301010b",
        1813 => x"67800000",
        1814 => x"93070004",
        1815 => x"232af900",
        1816 => x"93070002",
        1817 => x"a304f102",
        1818 => x"93070003",
        1819 => x"23220102",
        1820 => x"2305f102",
        1821 => x"23268100",
        1822 => x"930c5002",
        1823 => x"373b0000",
        1824 => x"b73b0000",
        1825 => x"373d0000",
        1826 => x"372c0000",
        1827 => x"930a0000",
        1828 => x"13840400",
        1829 => x"83470400",
        1830 => x"63840700",
        1831 => x"639c970d",
        1832 => x"b30d9440",
        1833 => x"63069402",
        1834 => x"93860d00",
        1835 => x"13860400",
        1836 => x"93050900",
        1837 => x"13050a00",
        1838 => x"eff01fbc",
        1839 => x"9307f0ff",
        1840 => x"6304f524",
        1841 => x"83274102",
        1842 => x"b387b701",
        1843 => x"2322f102",
        1844 => x"83470400",
        1845 => x"638a0722",
        1846 => x"9307f0ff",
        1847 => x"93041400",
        1848 => x"23280100",
        1849 => x"232e0100",
        1850 => x"232af100",
        1851 => x"232c0100",
        1852 => x"a3090104",
        1853 => x"23240106",
        1854 => x"930d1000",
        1855 => x"83c50400",
        1856 => x"13065000",
        1857 => x"13050be7",
        1858 => x"ef00d014",
        1859 => x"83270101",
        1860 => x"13841400",
        1861 => x"63140506",
        1862 => x"13f70701",
        1863 => x"63060700",
        1864 => x"13070002",
        1865 => x"a309e104",
        1866 => x"13f78700",
        1867 => x"63060700",
        1868 => x"1307b002",
        1869 => x"a309e104",
        1870 => x"83c60400",
        1871 => x"1307a002",
        1872 => x"638ce604",
        1873 => x"8327c101",
        1874 => x"13840400",
        1875 => x"93060000",
        1876 => x"13069000",
        1877 => x"1305a000",
        1878 => x"03470400",
        1879 => x"93051400",
        1880 => x"130707fd",
        1881 => x"637ee608",
        1882 => x"63840604",
        1883 => x"232ef100",
        1884 => x"6f000004",
        1885 => x"13041400",
        1886 => x"6ff0dff1",
        1887 => x"13070be7",
        1888 => x"3305e540",
        1889 => x"3395ad00",
        1890 => x"b3e7a700",
        1891 => x"2328f100",
        1892 => x"93040400",
        1893 => x"6ff09ff6",
        1894 => x"0327c100",
        1895 => x"93064700",
        1896 => x"03270700",
        1897 => x"2326d100",
        1898 => x"63420704",
        1899 => x"232ee100",
        1900 => x"03470400",
        1901 => x"9307e002",
        1902 => x"6314f708",
        1903 => x"03471400",
        1904 => x"9307a002",
        1905 => x"6318f704",
        1906 => x"8327c100",
        1907 => x"13042400",
        1908 => x"13874700",
        1909 => x"83a70700",
        1910 => x"2326e100",
        1911 => x"63d40700",
        1912 => x"9307f0ff",
        1913 => x"232af100",
        1914 => x"6f008005",
        1915 => x"3307e040",
        1916 => x"93e72700",
        1917 => x"232ee100",
        1918 => x"2328f100",
        1919 => x"6ff05ffb",
        1920 => x"b387a702",
        1921 => x"13840500",
        1922 => x"93061000",
        1923 => x"b387e700",
        1924 => x"6ff09ff4",
        1925 => x"13041400",
        1926 => x"232a0100",
        1927 => x"93060000",
        1928 => x"93070000",
        1929 => x"13069000",
        1930 => x"1305a000",
        1931 => x"03470400",
        1932 => x"93051400",
        1933 => x"130707fd",
        1934 => x"6372e608",
        1935 => x"e39406fa",
        1936 => x"83450400",
        1937 => x"13063000",
        1938 => x"13858be7",
        1939 => x"ef009000",
        1940 => x"63020502",
        1941 => x"93878be7",
        1942 => x"3305f540",
        1943 => x"83270101",
        1944 => x"13070004",
        1945 => x"3317a700",
        1946 => x"b3e7e700",
        1947 => x"13041400",
        1948 => x"2328f100",
        1949 => x"83450400",
        1950 => x"13066000",
        1951 => x"1305cde7",
        1952 => x"93041400",
        1953 => x"2304b102",
        1954 => x"ef00c07c",
        1955 => x"63080508",
        1956 => x"63980a04",
        1957 => x"03270101",
        1958 => x"8327c100",
        1959 => x"13770710",
        1960 => x"63080702",
        1961 => x"93874700",
        1962 => x"2326f100",
        1963 => x"83274102",
        1964 => x"b3873701",
        1965 => x"2322f102",
        1966 => x"6ff09fdd",
        1967 => x"b387a702",
        1968 => x"13840500",
        1969 => x"93061000",
        1970 => x"b387e700",
        1971 => x"6ff01ff6",
        1972 => x"93877700",
        1973 => x"93f787ff",
        1974 => x"93878700",
        1975 => x"6ff0dffc",
        1976 => x"1307c100",
        1977 => x"93068c87",
        1978 => x"13060900",
        1979 => x"93050101",
        1980 => x"13050a00",
        1981 => x"97000000",
        1982 => x"e7000000",
        1983 => x"9307f0ff",
        1984 => x"93090500",
        1985 => x"e314f5fa",
        1986 => x"8357c900",
        1987 => x"93f70704",
        1988 => x"e39407d0",
        1989 => x"03254102",
        1990 => x"6ff05fd0",
        1991 => x"1307c100",
        1992 => x"93068c87",
        1993 => x"13060900",
        1994 => x"93050101",
        1995 => x"13050a00",
        1996 => x"ef00801b",
        1997 => x"6ff09ffc",
        1998 => x"130101fd",
        1999 => x"232a5101",
        2000 => x"83a70501",
        2001 => x"930a0700",
        2002 => x"03a78500",
        2003 => x"23248102",
        2004 => x"23202103",
        2005 => x"232e3101",
        2006 => x"232c4101",
        2007 => x"23261102",
        2008 => x"23229102",
        2009 => x"23286101",
        2010 => x"23267101",
        2011 => x"93090500",
        2012 => x"13840500",
        2013 => x"13090600",
        2014 => x"138a0600",
        2015 => x"63d4e700",
        2016 => x"93070700",
        2017 => x"2320f900",
        2018 => x"03473404",
        2019 => x"63060700",
        2020 => x"93871700",
        2021 => x"2320f900",
        2022 => x"83270400",
        2023 => x"93f70702",
        2024 => x"63880700",
        2025 => x"83270900",
        2026 => x"93872700",
        2027 => x"2320f900",
        2028 => x"83240400",
        2029 => x"93f46400",
        2030 => x"639e0400",
        2031 => x"130b9401",
        2032 => x"930bf0ff",
        2033 => x"8327c400",
        2034 => x"03270900",
        2035 => x"b387e740",
        2036 => x"63c2f408",
        2037 => x"83473404",
        2038 => x"b336f000",
        2039 => x"83270400",
        2040 => x"93f70702",
        2041 => x"6390070c",
        2042 => x"13063404",
        2043 => x"93050a00",
        2044 => x"13850900",
        2045 => x"e7800a00",
        2046 => x"9307f0ff",
        2047 => x"6308f506",
        2048 => x"83270400",
        2049 => x"13074000",
        2050 => x"93040000",
        2051 => x"93f76700",
        2052 => x"639ce700",
        2053 => x"8324c400",
        2054 => x"83270900",
        2055 => x"b384f440",
        2056 => x"63d40400",
        2057 => x"93040000",
        2058 => x"83278400",
        2059 => x"03270401",
        2060 => x"6356f700",
        2061 => x"b387e740",
        2062 => x"b384f400",
        2063 => x"13090000",
        2064 => x"1304a401",
        2065 => x"130bf0ff",
        2066 => x"63902409",
        2067 => x"13050000",
        2068 => x"6f000002",
        2069 => x"93061000",
        2070 => x"13060b00",
        2071 => x"93050a00",
        2072 => x"13850900",
        2073 => x"e7800a00",
        2074 => x"631a7503",
        2075 => x"1305f0ff",
        2076 => x"8320c102",
        2077 => x"03248102",
        2078 => x"83244102",
        2079 => x"03290102",
        2080 => x"8329c101",
        2081 => x"032a8101",
        2082 => x"832a4101",
        2083 => x"032b0101",
        2084 => x"832bc100",
        2085 => x"13010103",
        2086 => x"67800000",
        2087 => x"93841400",
        2088 => x"6ff05ff2",
        2089 => x"3307d400",
        2090 => x"13060003",
        2091 => x"a301c704",
        2092 => x"03475404",
        2093 => x"93871600",
        2094 => x"b307f400",
        2095 => x"93862600",
        2096 => x"a381e704",
        2097 => x"6ff05ff2",
        2098 => x"93061000",
        2099 => x"13060400",
        2100 => x"93050a00",
        2101 => x"13850900",
        2102 => x"e7800a00",
        2103 => x"e30865f9",
        2104 => x"13091900",
        2105 => x"6ff05ff6",
        2106 => x"130101fd",
        2107 => x"23248102",
        2108 => x"23229102",
        2109 => x"23202103",
        2110 => x"232e3101",
        2111 => x"23261102",
        2112 => x"232c4101",
        2113 => x"232a5101",
        2114 => x"23286101",
        2115 => x"83c88501",
        2116 => x"93078007",
        2117 => x"93040500",
        2118 => x"13840500",
        2119 => x"13090600",
        2120 => x"93890600",
        2121 => x"63ee1701",
        2122 => x"93072006",
        2123 => x"93863504",
        2124 => x"63ee1701",
        2125 => x"638a082a",
        2126 => x"93078005",
        2127 => x"638af820",
        2128 => x"930a2404",
        2129 => x"23011405",
        2130 => x"6f004004",
        2131 => x"9387d8f9",
        2132 => x"93f7f70f",
        2133 => x"13065001",
        2134 => x"e364f6fe",
        2135 => x"37360000",
        2136 => x"93972700",
        2137 => x"1306c6ea",
        2138 => x"b387c700",
        2139 => x"83a70700",
        2140 => x"67800700",
        2141 => x"83270700",
        2142 => x"938a2504",
        2143 => x"93864700",
        2144 => x"83a70700",
        2145 => x"2320d700",
        2146 => x"2381f504",
        2147 => x"93071000",
        2148 => x"6f004029",
        2149 => x"03a60500",
        2150 => x"83270700",
        2151 => x"13750608",
        2152 => x"93854700",
        2153 => x"630e0504",
        2154 => x"83a70700",
        2155 => x"2320b700",
        2156 => x"37370000",
        2157 => x"83254400",
        2158 => x"130847e8",
        2159 => x"63d2071e",
        2160 => x"1307d002",
        2161 => x"a301e404",
        2162 => x"2324b400",
        2163 => x"63d80504",
        2164 => x"b307f040",
        2165 => x"1307a000",
        2166 => x"938a0600",
        2167 => x"33f6e702",
        2168 => x"938afaff",
        2169 => x"3306c800",
        2170 => x"03460600",
        2171 => x"2380ca00",
        2172 => x"13860700",
        2173 => x"b3d7e702",
        2174 => x"e372e6fe",
        2175 => x"6f008009",
        2176 => x"83a70700",
        2177 => x"13750604",
        2178 => x"2320b700",
        2179 => x"e30205fa",
        2180 => x"93970701",
        2181 => x"93d70741",
        2182 => x"6ff09ff9",
        2183 => x"1376b6ff",
        2184 => x"2320c400",
        2185 => x"6ff0dffa",
        2186 => x"03a60500",
        2187 => x"83270700",
        2188 => x"13750608",
        2189 => x"93854700",
        2190 => x"63080500",
        2191 => x"2320b700",
        2192 => x"83a70700",
        2193 => x"6f004001",
        2194 => x"13760604",
        2195 => x"2320b700",
        2196 => x"e30806fe",
        2197 => x"83d70700",
        2198 => x"37380000",
        2199 => x"1307f006",
        2200 => x"130848e8",
        2201 => x"639ae812",
        2202 => x"13078000",
        2203 => x"a3010404",
        2204 => x"03264400",
        2205 => x"2324c400",
        2206 => x"e34006f6",
        2207 => x"83250400",
        2208 => x"93f5b5ff",
        2209 => x"2320b400",
        2210 => x"e39807f4",
        2211 => x"938a0600",
        2212 => x"e31406f4",
        2213 => x"93078000",
        2214 => x"6314f702",
        2215 => x"83270400",
        2216 => x"93f71700",
        2217 => x"638e0700",
        2218 => x"03274400",
        2219 => x"83270401",
        2220 => x"63c8e700",
        2221 => x"93070003",
        2222 => x"a38ffafe",
        2223 => x"938afaff",
        2224 => x"b3865641",
        2225 => x"2328d400",
        2226 => x"13870900",
        2227 => x"93060900",
        2228 => x"1306c100",
        2229 => x"93050400",
        2230 => x"13850400",
        2231 => x"eff0dfc5",
        2232 => x"130af0ff",
        2233 => x"63164515",
        2234 => x"1305f0ff",
        2235 => x"8320c102",
        2236 => x"03248102",
        2237 => x"83244102",
        2238 => x"03290102",
        2239 => x"8329c101",
        2240 => x"032a8101",
        2241 => x"832a4101",
        2242 => x"032b0101",
        2243 => x"13010103",
        2244 => x"67800000",
        2245 => x"83a70500",
        2246 => x"93e70702",
        2247 => x"23a0f500",
        2248 => x"37380000",
        2249 => x"93088007",
        2250 => x"130888e9",
        2251 => x"03260400",
        2252 => x"a3021405",
        2253 => x"83270700",
        2254 => x"13750608",
        2255 => x"93854700",
        2256 => x"630e0500",
        2257 => x"2320b700",
        2258 => x"83a70700",
        2259 => x"6f000002",
        2260 => x"37380000",
        2261 => x"130848e8",
        2262 => x"6ff05ffd",
        2263 => x"13750604",
        2264 => x"2320b700",
        2265 => x"e30205fe",
        2266 => x"83d70700",
        2267 => x"13771600",
        2268 => x"63060700",
        2269 => x"13660602",
        2270 => x"2320c400",
        2271 => x"63860700",
        2272 => x"13070001",
        2273 => x"6ff09fee",
        2274 => x"03270400",
        2275 => x"1377f7fd",
        2276 => x"2320e400",
        2277 => x"6ff0dffe",
        2278 => x"1307a000",
        2279 => x"6ff01fed",
        2280 => x"130847e8",
        2281 => x"1307a000",
        2282 => x"6ff09fec",
        2283 => x"03a60500",
        2284 => x"83270700",
        2285 => x"83a54501",
        2286 => x"13780608",
        2287 => x"13854700",
        2288 => x"630a0800",
        2289 => x"2320a700",
        2290 => x"83a70700",
        2291 => x"23a0b700",
        2292 => x"6f008001",
        2293 => x"2320a700",
        2294 => x"13760604",
        2295 => x"83a70700",
        2296 => x"e30606fe",
        2297 => x"2390b700",
        2298 => x"23280400",
        2299 => x"938a0600",
        2300 => x"6ff09fed",
        2301 => x"83270700",
        2302 => x"03a64500",
        2303 => x"93050000",
        2304 => x"93864700",
        2305 => x"2320d700",
        2306 => x"83aa0700",
        2307 => x"13850a00",
        2308 => x"ef004024",
        2309 => x"63060500",
        2310 => x"33055541",
        2311 => x"2322a400",
        2312 => x"83274400",
        2313 => x"2328f400",
        2314 => x"a3010404",
        2315 => x"6ff0dfe9",
        2316 => x"83260401",
        2317 => x"13860a00",
        2318 => x"93050900",
        2319 => x"13850400",
        2320 => x"e7800900",
        2321 => x"e30245eb",
        2322 => x"83270400",
        2323 => x"93f72700",
        2324 => x"63940704",
        2325 => x"8327c100",
        2326 => x"0325c400",
        2327 => x"e358f5e8",
        2328 => x"13850700",
        2329 => x"6ff09fe8",
        2330 => x"93061000",
        2331 => x"13860a00",
        2332 => x"93050900",
        2333 => x"13850400",
        2334 => x"e7800900",
        2335 => x"e30665e7",
        2336 => x"130a1a00",
        2337 => x"8327c400",
        2338 => x"0327c100",
        2339 => x"b387e740",
        2340 => x"e34cfafc",
        2341 => x"6ff01ffc",
        2342 => x"130a0000",
        2343 => x"930a9401",
        2344 => x"130bf0ff",
        2345 => x"6ff01ffe",
        2346 => x"130101ff",
        2347 => x"23248100",
        2348 => x"13840500",
        2349 => x"83a50500",
        2350 => x"23229100",
        2351 => x"23261100",
        2352 => x"93040500",
        2353 => x"63840500",
        2354 => x"eff01ffe",
        2355 => x"93050400",
        2356 => x"03248100",
        2357 => x"8320c100",
        2358 => x"13850400",
        2359 => x"83244100",
        2360 => x"13010101",
        2361 => x"6f004019",
        2362 => x"83a7c187",
        2363 => x"6382a716",
        2364 => x"83274502",
        2365 => x"130101fe",
        2366 => x"232c8100",
        2367 => x"232e1100",
        2368 => x"232a9100",
        2369 => x"23282101",
        2370 => x"23263101",
        2371 => x"13040500",
        2372 => x"638a0704",
        2373 => x"83a7c700",
        2374 => x"638c0702",
        2375 => x"93040000",
        2376 => x"13090008",
        2377 => x"83274402",
        2378 => x"83a7c700",
        2379 => x"b3879700",
        2380 => x"83a50700",
        2381 => x"6396050e",
        2382 => x"93844400",
        2383 => x"e39424ff",
        2384 => x"83274402",
        2385 => x"13050400",
        2386 => x"83a5c700",
        2387 => x"ef00c012",
        2388 => x"83274402",
        2389 => x"83a50700",
        2390 => x"63860500",
        2391 => x"13050400",
        2392 => x"ef008011",
        2393 => x"83254401",
        2394 => x"63860500",
        2395 => x"13050400",
        2396 => x"ef008010",
        2397 => x"83254402",
        2398 => x"63860500",
        2399 => x"13050400",
        2400 => x"ef00800f",
        2401 => x"83258403",
        2402 => x"63860500",
        2403 => x"13050400",
        2404 => x"ef00800e",
        2405 => x"8325c403",
        2406 => x"63860500",
        2407 => x"13050400",
        2408 => x"ef00800d",
        2409 => x"83250404",
        2410 => x"63860500",
        2411 => x"13050400",
        2412 => x"ef00800c",
        2413 => x"8325c405",
        2414 => x"63860500",
        2415 => x"13050400",
        2416 => x"ef00800b",
        2417 => x"83258405",
        2418 => x"63860500",
        2419 => x"13050400",
        2420 => x"ef00800a",
        2421 => x"83254403",
        2422 => x"63860500",
        2423 => x"13050400",
        2424 => x"ef008009",
        2425 => x"83278401",
        2426 => x"63860704",
        2427 => x"83278402",
        2428 => x"13050400",
        2429 => x"e7800700",
        2430 => x"83258404",
        2431 => x"638c0502",
        2432 => x"13050400",
        2433 => x"03248101",
        2434 => x"8320c101",
        2435 => x"83244101",
        2436 => x"03290101",
        2437 => x"8329c100",
        2438 => x"13010102",
        2439 => x"6ff0dfe8",
        2440 => x"83a90500",
        2441 => x"13050400",
        2442 => x"ef000005",
        2443 => x"93850900",
        2444 => x"6ff05ff0",
        2445 => x"8320c101",
        2446 => x"03248101",
        2447 => x"83244101",
        2448 => x"03290101",
        2449 => x"8329c100",
        2450 => x"13010102",
        2451 => x"67800000",
        2452 => x"67800000",
        2453 => x"93f5f50f",
        2454 => x"3306c500",
        2455 => x"6316c500",
        2456 => x"13050000",
        2457 => x"67800000",
        2458 => x"83470500",
        2459 => x"e38cb7fe",
        2460 => x"13051500",
        2461 => x"6ff09ffe",
        2462 => x"638a050e",
        2463 => x"83a7c5ff",
        2464 => x"130101fe",
        2465 => x"232c8100",
        2466 => x"232e1100",
        2467 => x"1384c5ff",
        2468 => x"63d40700",
        2469 => x"3304f400",
        2470 => x"2326a100",
        2471 => x"ef008033",
        2472 => x"83a7c188",
        2473 => x"0325c100",
        2474 => x"639e0700",
        2475 => x"23220400",
        2476 => x"23a68188",
        2477 => x"03248101",
        2478 => x"8320c101",
        2479 => x"13010102",
        2480 => x"6f008031",
        2481 => x"6374f402",
        2482 => x"03260400",
        2483 => x"b306c400",
        2484 => x"639ad700",
        2485 => x"83a60700",
        2486 => x"83a74700",
        2487 => x"b386c600",
        2488 => x"2320d400",
        2489 => x"2322f400",
        2490 => x"6ff09ffc",
        2491 => x"13870700",
        2492 => x"83a74700",
        2493 => x"63840700",
        2494 => x"e37af4fe",
        2495 => x"83260700",
        2496 => x"3306d700",
        2497 => x"63188602",
        2498 => x"03260400",
        2499 => x"b386c600",
        2500 => x"2320d700",
        2501 => x"3306d700",
        2502 => x"e39ec7f8",
        2503 => x"03a60700",
        2504 => x"83a74700",
        2505 => x"b306d600",
        2506 => x"2320d700",
        2507 => x"2322f700",
        2508 => x"6ff05ff8",
        2509 => x"6378c400",
        2510 => x"9307c000",
        2511 => x"2320f500",
        2512 => x"6ff05ff7",
        2513 => x"03260400",
        2514 => x"b306c400",
        2515 => x"639ad700",
        2516 => x"83a60700",
        2517 => x"83a74700",
        2518 => x"b386c600",
        2519 => x"2320d400",
        2520 => x"2322f400",
        2521 => x"23228700",
        2522 => x"6ff0dff4",
        2523 => x"67800000",
        2524 => x"130101fe",
        2525 => x"232a9100",
        2526 => x"93843500",
        2527 => x"93f4c4ff",
        2528 => x"23282101",
        2529 => x"232e1100",
        2530 => x"232c8100",
        2531 => x"23263101",
        2532 => x"93848400",
        2533 => x"9307c000",
        2534 => x"13090500",
        2535 => x"63f0f406",
        2536 => x"9304c000",
        2537 => x"63eeb404",
        2538 => x"13050900",
        2539 => x"ef008022",
        2540 => x"03a7c188",
        2541 => x"13040700",
        2542 => x"63180406",
        2543 => x"83a78188",
        2544 => x"639a0700",
        2545 => x"93050000",
        2546 => x"13050900",
        2547 => x"ef00001c",
        2548 => x"23a4a188",
        2549 => x"93850400",
        2550 => x"13050900",
        2551 => x"ef00001b",
        2552 => x"9309f0ff",
        2553 => x"631a350b",
        2554 => x"9307c000",
        2555 => x"2320f900",
        2556 => x"13050900",
        2557 => x"ef00401e",
        2558 => x"6f000001",
        2559 => x"e3d404fa",
        2560 => x"9307c000",
        2561 => x"2320f900",
        2562 => x"13050000",
        2563 => x"8320c101",
        2564 => x"03248101",
        2565 => x"83244101",
        2566 => x"03290101",
        2567 => x"8329c100",
        2568 => x"13010102",
        2569 => x"67800000",
        2570 => x"83270400",
        2571 => x"b3879740",
        2572 => x"63ce0704",
        2573 => x"1306b000",
        2574 => x"637af600",
        2575 => x"2320f400",
        2576 => x"3304f400",
        2577 => x"23209400",
        2578 => x"6f000001",
        2579 => x"83274400",
        2580 => x"631a8702",
        2581 => x"23a6f188",
        2582 => x"13050900",
        2583 => x"ef00c017",
        2584 => x"1305b400",
        2585 => x"93074400",
        2586 => x"137585ff",
        2587 => x"3307f540",
        2588 => x"e30ef5f8",
        2589 => x"3304e400",
        2590 => x"b387a740",
        2591 => x"2320f400",
        2592 => x"6ff0dff8",
        2593 => x"2322f700",
        2594 => x"6ff01ffd",
        2595 => x"13070400",
        2596 => x"03244400",
        2597 => x"6ff05ff2",
        2598 => x"13043500",
        2599 => x"1374c4ff",
        2600 => x"e30285fa",
        2601 => x"b305a440",
        2602 => x"13050900",
        2603 => x"ef00000e",
        2604 => x"e31a35f9",
        2605 => x"6ff05ff3",
        2606 => x"130101fe",
        2607 => x"232c8100",
        2608 => x"232e1100",
        2609 => x"232a9100",
        2610 => x"23282101",
        2611 => x"23263101",
        2612 => x"23244101",
        2613 => x"13040600",
        2614 => x"63940502",
        2615 => x"03248101",
        2616 => x"8320c101",
        2617 => x"83244101",
        2618 => x"03290101",
        2619 => x"8329c100",
        2620 => x"032a8100",
        2621 => x"93050600",
        2622 => x"13010102",
        2623 => x"6ff05fe7",
        2624 => x"63180602",
        2625 => x"eff05fd7",
        2626 => x"93040000",
        2627 => x"8320c101",
        2628 => x"03248101",
        2629 => x"03290101",
        2630 => x"8329c100",
        2631 => x"032a8100",
        2632 => x"13850400",
        2633 => x"83244101",
        2634 => x"13010102",
        2635 => x"67800000",
        2636 => x"130a0500",
        2637 => x"93840500",
        2638 => x"ef00400a",
        2639 => x"13090500",
        2640 => x"63668500",
        2641 => x"93571500",
        2642 => x"e3e287fc",
        2643 => x"93050400",
        2644 => x"13050a00",
        2645 => x"eff0dfe1",
        2646 => x"93090500",
        2647 => x"e30605fa",
        2648 => x"13060400",
        2649 => x"63748900",
        2650 => x"13060900",
        2651 => x"93850400",
        2652 => x"13850900",
        2653 => x"efe05f97",
        2654 => x"93850400",
        2655 => x"13050a00",
        2656 => x"eff09fcf",
        2657 => x"93840900",
        2658 => x"6ff05ff8",
        2659 => x"130101ff",
        2660 => x"23248100",
        2661 => x"23229100",
        2662 => x"13040500",
        2663 => x"13850500",
        2664 => x"23261100",
        2665 => x"23a20188",
        2666 => x"ef00000c",
        2667 => x"9307f0ff",
        2668 => x"6318f500",
        2669 => x"83a74188",
        2670 => x"63840700",
        2671 => x"2320f400",
        2672 => x"8320c100",
        2673 => x"03248100",
        2674 => x"83244100",
        2675 => x"13010101",
        2676 => x"67800000",
        2677 => x"67800000",
        2678 => x"67800000",
        2679 => x"83a7c5ff",
        2680 => x"1385c7ff",
        2681 => x"63d80700",
        2682 => x"b385a500",
        2683 => x"83a70500",
        2684 => x"3305f500",
        2685 => x"67800000",
        2686 => x"9308d005",
        2687 => x"73000000",
        2688 => x"63520502",
        2689 => x"130101ff",
        2690 => x"23248100",
        2691 => x"13040500",
        2692 => x"23261100",
        2693 => x"33048040",
        2694 => x"efe0dfc4",
        2695 => x"23208500",
        2696 => x"6f000000",
        2697 => x"6f000000",
        2698 => x"130101ff",
        2699 => x"23261100",
        2700 => x"23248100",
        2701 => x"9308900a",
        2702 => x"73000000",
        2703 => x"13040500",
        2704 => x"635a0500",
        2705 => x"33048040",
        2706 => x"efe0dfc1",
        2707 => x"23208500",
        2708 => x"1304f0ff",
        2709 => x"8320c100",
        2710 => x"13050400",
        2711 => x"03248100",
        2712 => x"13010101",
        2713 => x"67800000",
        2714 => x"03a70189",
        2715 => x"130101ff",
        2716 => x"23261100",
        2717 => x"93070500",
        2718 => x"631c0702",
        2719 => x"9308600d",
        2720 => x"13050000",
        2721 => x"73000000",
        2722 => x"1307f0ff",
        2723 => x"6310e502",
        2724 => x"efe05fbd",
        2725 => x"9307c000",
        2726 => x"2320f500",
        2727 => x"1305f0ff",
        2728 => x"8320c100",
        2729 => x"13010101",
        2730 => x"67800000",
        2731 => x"23a8a188",
        2732 => x"03a70189",
        2733 => x"9308600d",
        2734 => x"b387e700",
        2735 => x"13850700",
        2736 => x"73000000",
        2737 => x"e316f5fc",
        2738 => x"23a8a188",
        2739 => x"13050700",
        2740 => x"6ff01ffd",
        2741 => x"10000000",
        2742 => x"00000000",
        2743 => x"037a5200",
        2744 => x"017c0101",
        2745 => x"1b0d0200",
        2746 => x"10000000",
        2747 => x"18000000",
        2748 => x"6cdbffff",
        2749 => x"78040000",
        2750 => x"00000000",
        2751 => x"10000000",
        2752 => x"00000000",
        2753 => x"037a5200",
        2754 => x"017c0101",
        2755 => x"1b0d0200",
        2756 => x"10000000",
        2757 => x"18000000",
        2758 => x"bcdfffff",
        2759 => x"30040000",
        2760 => x"00000000",
        2761 => x"10000000",
        2762 => x"00000000",
        2763 => x"037a5200",
        2764 => x"017c0101",
        2765 => x"1b0d0200",
        2766 => x"10000000",
        2767 => x"18000000",
        2768 => x"c4e3ffff",
        2769 => x"e4030000",
        2770 => x"00000000",
        2771 => x"c0030000",
        2772 => x"9c030000",
        2773 => x"b4030000",
        2774 => x"a8030000",
        2775 => x"f0020000",
        2776 => x"f0020000",
        2777 => x"f0020000",
        2778 => x"04040000",
        2779 => x"f0020000",
        2780 => x"f0020000",
        2781 => x"f0020000",
        2782 => x"f0020000",
        2783 => x"f0020000",
        2784 => x"f0020000",
        2785 => x"f0020000",
        2786 => x"cc030000",
        2787 => x"68040000",
        2788 => x"20040000",
        2789 => x"20040000",
        2790 => x"20040000",
        2791 => x"20040000",
        2792 => x"5c040000",
        2793 => x"a8040000",
        2794 => x"80040000",
        2795 => x"20040000",
        2796 => x"20040000",
        2797 => x"20040000",
        2798 => x"20040000",
        2799 => x"20040000",
        2800 => x"20040000",
        2801 => x"20040000",
        2802 => x"20040000",
        2803 => x"20040000",
        2804 => x"20040000",
        2805 => x"20040000",
        2806 => x"20040000",
        2807 => x"20040000",
        2808 => x"20040000",
        2809 => x"48040000",
        2810 => x"48040000",
        2811 => x"20040000",
        2812 => x"20040000",
        2813 => x"20040000",
        2814 => x"20040000",
        2815 => x"20040000",
        2816 => x"20040000",
        2817 => x"20040000",
        2818 => x"20040000",
        2819 => x"20040000",
        2820 => x"20040000",
        2821 => x"20040000",
        2822 => x"20040000",
        2823 => x"5c040000",
        2824 => x"68040000",
        2825 => x"24050000",
        2826 => x"0c050000",
        2827 => x"20040000",
        2828 => x"20040000",
        2829 => x"20040000",
        2830 => x"20040000",
        2831 => x"20040000",
        2832 => x"20040000",
        2833 => x"f4040000",
        2834 => x"20040000",
        2835 => x"20040000",
        2836 => x"20040000",
        2837 => x"20040000",
        2838 => x"48040000",
        2839 => x"48040000",
        2840 => x"00010202",
        2841 => x"03030303",
        2842 => x"04040404",
        2843 => x"04040404",
        2844 => x"05050505",
        2845 => x"05050505",
        2846 => x"05050505",
        2847 => x"05050505",
        2848 => x"06060606",
        2849 => x"06060606",
        2850 => x"06060606",
        2851 => x"06060606",
        2852 => x"06060606",
        2853 => x"06060606",
        2854 => x"06060606",
        2855 => x"06060606",
        2856 => x"07070707",
        2857 => x"07070707",
        2858 => x"07070707",
        2859 => x"07070707",
        2860 => x"07070707",
        2861 => x"07070707",
        2862 => x"07070707",
        2863 => x"07070707",
        2864 => x"07070707",
        2865 => x"07070707",
        2866 => x"07070707",
        2867 => x"07070707",
        2868 => x"07070707",
        2869 => x"07070707",
        2870 => x"07070707",
        2871 => x"07070707",
        2872 => x"08080808",
        2873 => x"08080808",
        2874 => x"08080808",
        2875 => x"08080808",
        2876 => x"08080808",
        2877 => x"08080808",
        2878 => x"08080808",
        2879 => x"08080808",
        2880 => x"08080808",
        2881 => x"08080808",
        2882 => x"08080808",
        2883 => x"08080808",
        2884 => x"08080808",
        2885 => x"08080808",
        2886 => x"08080808",
        2887 => x"08080808",
        2888 => x"08080808",
        2889 => x"08080808",
        2890 => x"08080808",
        2891 => x"08080808",
        2892 => x"08080808",
        2893 => x"08080808",
        2894 => x"08080808",
        2895 => x"08080808",
        2896 => x"08080808",
        2897 => x"08080808",
        2898 => x"08080808",
        2899 => x"08080808",
        2900 => x"08080808",
        2901 => x"08080808",
        2902 => x"08080808",
        2903 => x"08080808",
        2904 => x"0d0a4542",
        2905 => x"5245414b",
        2906 => x"21206d69",
        2907 => x"70203d20",
        2908 => x"00000000",
        2909 => x"0d0a0d0a",
        2910 => x"44697370",
        2911 => x"6c617969",
        2912 => x"6e672074",
        2913 => x"68652074",
        2914 => x"696d6520",
        2915 => x"70617373",
        2916 => x"65642073",
        2917 => x"696e6365",
        2918 => x"20726573",
        2919 => x"65740d0a",
        2920 => x"0d0a0000",
        2921 => x"2530356c",
        2922 => x"643a2530",
        2923 => x"366c6420",
        2924 => x"20202530",
        2925 => x"326c643a",
        2926 => x"2530326c",
        2927 => x"643a2530",
        2928 => x"326c640d",
        2929 => x"00000000",
        2930 => x"696e7465",
        2931 => x"72727570",
        2932 => x"745f6469",
        2933 => x"72656374",
        2934 => x"00000000",
        2935 => x"54485541",
        2936 => x"53205249",
        2937 => x"53432d56",
        2938 => x"20525633",
        2939 => x"32494d20",
        2940 => x"62617265",
        2941 => x"206d6574",
        2942 => x"616c2070",
        2943 => x"726f6365",
        2944 => x"73736f72",
        2945 => x"00000000",
        2946 => x"54686520",
        2947 => x"48616775",
        2948 => x"6520556e",
        2949 => x"69766572",
        2950 => x"73697479",
        2951 => x"206f6620",
        2952 => x"4170706c",
        2953 => x"69656420",
        2954 => x"53636965",
        2955 => x"6e636573",
        2956 => x"00000000",
        2957 => x"44657061",
        2958 => x"72746d65",
        2959 => x"6e74206f",
        2960 => x"6620456c",
        2961 => x"65637472",
        2962 => x"6963616c",
        2963 => x"20456e67",
        2964 => x"696e6565",
        2965 => x"72696e67",
        2966 => x"00000000",
        2967 => x"4a2e452e",
        2968 => x"4a2e206f",
        2969 => x"70206465",
        2970 => x"6e204272",
        2971 => x"6f757700",
        2972 => x"232d302b",
        2973 => x"20000000",
        2974 => x"686c4c00",
        2975 => x"65666745",
        2976 => x"46470000",
        2977 => x"30313233",
        2978 => x"34353637",
        2979 => x"38394142",
        2980 => x"43444546",
        2981 => x"00000000",
        2982 => x"30313233",
        2983 => x"34353637",
        2984 => x"38396162",
        2985 => x"63646566",
        2986 => x"00000000",
        2987 => x"74210000",
        2988 => x"94210000",
        2989 => x"40210000",
        2990 => x"40210000",
        2991 => x"40210000",
        2992 => x"40210000",
        2993 => x"94210000",
        2994 => x"40210000",
        2995 => x"40210000",
        2996 => x"40210000",
        2997 => x"40210000",
        2998 => x"ac230000",
        2999 => x"28220000",
        3000 => x"14230000",
        3001 => x"40210000",
        3002 => x"40210000",
        3003 => x"f4230000",
        3004 => x"40210000",
        3005 => x"28220000",
        3006 => x"40210000",
        3007 => x"40210000",
        3008 => x"20230000",
        3009 => x"18000020",
        3010 => x"c82d0000",
        3011 => x"dc2d0000",
        3012 => x"082e0000",
        3013 => x"342e0000",
        3014 => x"5c2e0000",
        3015 => x"00000000",
        3016 => x"00000000",
        3017 => x"00000000",
        3018 => x"00000000",
        3019 => x"00000000",
        3020 => x"00000000",
        3021 => x"00000000",
        3022 => x"00000000",
        3023 => x"00000000",
        3024 => x"00000000",
        3025 => x"00000000",
        3026 => x"00000000",
        3027 => x"00000000",
        3028 => x"00000000",
        3029 => x"00000000",
        3030 => x"00000000",
        3031 => x"00000000",
        3032 => x"00000000",
        3033 => x"00000000",
        3034 => x"00000000",
        3035 => x"00000000",
        3036 => x"00000000",
        3037 => x"00000000",
        3038 => x"00000000",
        3039 => x"00000000",
        3040 => x"80000020",
        3041 => x"18000020",
        others => (others => '0')
    );
end package processor_common_rom;
