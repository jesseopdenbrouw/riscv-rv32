-- #################################################################################################
-- # bootloader.vhd - The bootloader ROM                                                           #
-- # ********************************************************************************************* #
-- # This file is part of the THUAS RISCV RV32 Project                                             #
-- # ********************************************************************************************* #
-- # BSD 3-Clause License                                                                          #
-- #                                                                                               #
-- # Copyright (c) 2023, Jesse op den Brouw. All rights reserved.                                  #
-- #                                                                                               #
-- # Redistribution and use in source and binary forms, with or without modification, are          #
-- # permitted provided that the following conditions are met:                                     #
-- #                                                                                               #
-- # 1. Redistributions of source code must retain the above copyright notice, this list of        #
-- #    conditions and the following disclaimer.                                                   #
-- #                                                                                               #
-- # 2. Redistributions in binary form must reproduce the above copyright notice, this list of     #
-- #    conditions and the following disclaimer in the documentation and/or other materials        #
-- #    provided with the distribution.                                                            #
-- #                                                                                               #
-- # 3. Neither the name of the copyright holder nor the names of its contributors may be used to  #
-- #    endorse or promote products derived from this software without specific prior written      #
-- #    permission.                                                                                #
-- #                                                                                               #
-- # THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND ANY EXPRESS   #
-- # OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED WARRANTIES OF               #
-- # MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE    #
-- # COPYRIGHT HOLDER OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL,     #
-- # EXEMPLARY, OR CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE #
-- # GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER CAUSED    #
-- # AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT (INCLUDING     #
-- # NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED  #
-- # OF THE POSSIBILITY OF SUCH DAMAGE.                                                            #
-- # ********************************************************************************************* #
-- # https:/github.com/jesseopdenbrouw/riscv-rv32                                                  #
-- #################################################################################################

-- This file contains the description of the bootloader ROM. The ROM
-- is placed in immutable onboard RAM blocks. A read takes two
-- clock cycles, for both instruction and data.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.processor_common.all;
use work.processor_common_rom.all;

entity bootloader is
    port (I_clk : in std_logic;
          I_areset : in std_logic;
          I_pc : in data_type;
          I_memaddress : in data_type;
          I_memsize : in memsize_type;
          I_csboot : in std_logic;
          I_stall : in std_logic;
          O_instr : out data_type;
          O_dataout : out data_type;
          --
          O_load_misaligned_error : out std_logic
         );
end entity bootloader;

architecture rtl of bootloader is

-- The bootloader ROM
signal bootrom : bootloader_type := (
           0 => x"97020000",
           1 => x"9382c207",
           2 => x"73905230",
           3 => x"97010010",
           4 => x"9381417f",
           5 => x"17810010",
           6 => x"1301c1fe",
           7 => x"93878186",
           8 => x"13874186",
           9 => x"13060000",
          10 => x"63e4e700",
          11 => x"3386e740",
          12 => x"93050000",
          13 => x"13854186",
          14 => x"ef00c006",
          15 => x"37050020",
          16 => x"93874186",
          17 => x"13070500",
          18 => x"13060000",
          19 => x"63e4e700",
          20 => x"3386e740",
          21 => x"b7150010",
          22 => x"938585e7",
          23 => x"13050500",
          24 => x"ef000002",
          25 => x"ef00d025",
          26 => x"13060000",
          27 => x"93854186",
          28 => x"13050000",
          29 => x"ef00c051",
          30 => x"ef009020",
          31 => x"6f000000",
          32 => x"13030500",
          33 => x"630e0600",
          34 => x"83830500",
          35 => x"23007300",
          36 => x"1306f6ff",
          37 => x"13031300",
          38 => x"93851500",
          39 => x"e31606fe",
          40 => x"67800000",
          41 => x"13030500",
          42 => x"630a0600",
          43 => x"2300b300",
          44 => x"1306f6ff",
          45 => x"13031300",
          46 => x"e31a06fe",
          47 => x"67800000",
          48 => x"03460500",
          49 => x"83c60500",
          50 => x"13051500",
          51 => x"93851500",
          52 => x"6314d600",
          53 => x"e31606fe",
          54 => x"3305d640",
          55 => x"67800000",
          56 => x"6f000000",
          57 => x"b70700f0",
          58 => x"03a54702",
          59 => x"13754500",
          60 => x"67800000",
          61 => x"370700f0",
          62 => x"83274702",
          63 => x"93f74700",
          64 => x"e38c07fe",
          65 => x"03258702",
          66 => x"1375f50f",
          67 => x"67800000",
          68 => x"130101fd",
          69 => x"23202103",
          70 => x"37190010",
          71 => x"23248102",
          72 => x"23229102",
          73 => x"232e3101",
          74 => x"232c4101",
          75 => x"232a5101",
          76 => x"23286101",
          77 => x"23267101",
          78 => x"23248101",
          79 => x"23261102",
          80 => x"93040500",
          81 => x"13040000",
          82 => x"130949bb",
          83 => x"930a5001",
          84 => x"938bf5ff",
          85 => x"130bf007",
          86 => x"130a2000",
          87 => x"93092001",
          88 => x"371c0010",
          89 => x"eff01ff9",
          90 => x"1377f50f",
          91 => x"63c4ea0a",
          92 => x"6354ea04",
          93 => x"9307d7ff",
          94 => x"63e0f904",
          95 => x"93972700",
          96 => x"b307f900",
          97 => x"83a70700",
          98 => x"67800700",
          99 => x"630a0400",
         100 => x"1304f4ff",
         101 => x"1305f007",
         102 => x"ef000013",
         103 => x"e31a04fe",
         104 => x"eff05ff5",
         105 => x"1377f50f",
         106 => x"13040000",
         107 => x"e3d2eafc",
         108 => x"9307f007",
         109 => x"630ef70c",
         110 => x"63547405",
         111 => x"9377f50f",
         112 => x"938607fe",
         113 => x"93f6f60f",
         114 => x"1306e005",
         115 => x"e36cd6f8",
         116 => x"b3868400",
         117 => x"13050700",
         118 => x"2380f600",
         119 => x"ef00c00e",
         120 => x"eff05ff1",
         121 => x"1377f50f",
         122 => x"93075001",
         123 => x"13041400",
         124 => x"e3d0e7f8",
         125 => x"9307f007",
         126 => x"6302f702",
         127 => x"e34074fd",
         128 => x"13057000",
         129 => x"ef00400c",
         130 => x"eff0dfee",
         131 => x"1377f50f",
         132 => x"e3d0eaf6",
         133 => x"e31267fb",
         134 => x"630c0406",
         135 => x"1305f007",
         136 => x"ef00800a",
         137 => x"1304f4ff",
         138 => x"6ff0dff3",
         139 => x"b3848400",
         140 => x"37150010",
         141 => x"23800400",
         142 => x"130505c2",
         143 => x"ef00c00a",
         144 => x"8320c102",
         145 => x"13050400",
         146 => x"03248102",
         147 => x"83244102",
         148 => x"03290102",
         149 => x"8329c101",
         150 => x"032a8101",
         151 => x"832a4101",
         152 => x"032b0101",
         153 => x"832bc100",
         154 => x"032c8100",
         155 => x"13010103",
         156 => x"67800000",
         157 => x"13058ce6",
         158 => x"ef000007",
         159 => x"eff09fe7",
         160 => x"1377f50f",
         161 => x"13040000",
         162 => x"e3d4eaee",
         163 => x"6ff05ff2",
         164 => x"13057000",
         165 => x"ef004003",
         166 => x"6ff09ff0",
         167 => x"f32710fc",
         168 => x"63960700",
         169 => x"b7f7fa02",
         170 => x"93870708",
         171 => x"63060500",
         172 => x"33d5a702",
         173 => x"1305f5ff",
         174 => x"b70700f0",
         175 => x"23a6a702",
         176 => x"23a0b702",
         177 => x"67800000",
         178 => x"1375f50f",
         179 => x"b70700f0",
         180 => x"370700f0",
         181 => x"23a4a702",
         182 => x"83274702",
         183 => x"93f70701",
         184 => x"e38c07fe",
         185 => x"67800000",
         186 => x"630e0502",
         187 => x"130101ff",
         188 => x"23248100",
         189 => x"23261100",
         190 => x"13040500",
         191 => x"03450500",
         192 => x"630a0500",
         193 => x"13041400",
         194 => x"eff01ffc",
         195 => x"03450400",
         196 => x"e31a05fe",
         197 => x"8320c100",
         198 => x"03248100",
         199 => x"13010101",
         200 => x"67800000",
         201 => x"67800000",
         202 => x"130101fe",
         203 => x"232e1100",
         204 => x"232c8100",
         205 => x"232a9100",
         206 => x"23282101",
         207 => x"23263101",
         208 => x"23244101",
         209 => x"6358a008",
         210 => x"b7190010",
         211 => x"13090500",
         212 => x"93040000",
         213 => x"13040000",
         214 => x"938959d6",
         215 => x"130a1000",
         216 => x"6f000001",
         217 => x"3364c400",
         218 => x"93841400",
         219 => x"63029904",
         220 => x"eff05fd8",
         221 => x"b387a900",
         222 => x"83c70700",
         223 => x"130605fd",
         224 => x"13144400",
         225 => x"13f74700",
         226 => x"93f64704",
         227 => x"e31c07fc",
         228 => x"93f73700",
         229 => x"e38a06fc",
         230 => x"63944701",
         231 => x"13050502",
         232 => x"130595fa",
         233 => x"93841400",
         234 => x"3364a400",
         235 => x"e31299fc",
         236 => x"8320c101",
         237 => x"13050400",
         238 => x"03248101",
         239 => x"83244101",
         240 => x"03290101",
         241 => x"8329c100",
         242 => x"032a8100",
         243 => x"13010102",
         244 => x"67800000",
         245 => x"13040000",
         246 => x"6ff09ffd",
         247 => x"83470500",
         248 => x"37160010",
         249 => x"130656d6",
         250 => x"3307f600",
         251 => x"03470700",
         252 => x"93060500",
         253 => x"13758700",
         254 => x"630e0500",
         255 => x"83c71600",
         256 => x"93861600",
         257 => x"3307f600",
         258 => x"03470700",
         259 => x"13758700",
         260 => x"e31605fe",
         261 => x"13754704",
         262 => x"630a0506",
         263 => x"13050000",
         264 => x"13031000",
         265 => x"6f000002",
         266 => x"83c71600",
         267 => x"33e5a800",
         268 => x"93861600",
         269 => x"3307f600",
         270 => x"03470700",
         271 => x"13784704",
         272 => x"63000804",
         273 => x"13784700",
         274 => x"938807fd",
         275 => x"13773700",
         276 => x"13154500",
         277 => x"e31a08fc",
         278 => x"63146700",
         279 => x"93870702",
         280 => x"938797fa",
         281 => x"33e5a700",
         282 => x"83c71600",
         283 => x"93861600",
         284 => x"3307f600",
         285 => x"03470700",
         286 => x"13784704",
         287 => x"e31408fc",
         288 => x"63840500",
         289 => x"23a0d500",
         290 => x"67800000",
         291 => x"13050000",
         292 => x"6ff01fff",
         293 => x"130101fe",
         294 => x"232e1100",
         295 => x"232c8100",
         296 => x"23220100",
         297 => x"23240100",
         298 => x"23260100",
         299 => x"63000506",
         300 => x"13040500",
         301 => x"63440504",
         302 => x"93074100",
         303 => x"9306a000",
         304 => x"93059000",
         305 => x"3377d402",
         306 => x"13850700",
         307 => x"9387f7ff",
         308 => x"13060400",
         309 => x"13070703",
         310 => x"a385e700",
         311 => x"3354d402",
         312 => x"e3e2c5fe",
         313 => x"3305d500",
         314 => x"eff01fe0",
         315 => x"8320c101",
         316 => x"03248101",
         317 => x"13010102",
         318 => x"67800000",
         319 => x"1305d002",
         320 => x"eff09fdc",
         321 => x"33048040",
         322 => x"6ff01ffb",
         323 => x"13050003",
         324 => x"eff09fdb",
         325 => x"8320c101",
         326 => x"03248101",
         327 => x"13010102",
         328 => x"67800000",
         329 => x"130101fe",
         330 => x"232e1100",
         331 => x"23220100",
         332 => x"23240100",
         333 => x"23060100",
         334 => x"9387f5ff",
         335 => x"13077000",
         336 => x"6376f700",
         337 => x"93077000",
         338 => x"93058000",
         339 => x"13074100",
         340 => x"b307f700",
         341 => x"b385b740",
         342 => x"13069003",
         343 => x"9376f500",
         344 => x"13870603",
         345 => x"6374e600",
         346 => x"13877605",
         347 => x"2380e700",
         348 => x"9387f7ff",
         349 => x"13554500",
         350 => x"e392f5fe",
         351 => x"13054100",
         352 => x"eff09fd6",
         353 => x"8320c101",
         354 => x"13010102",
         355 => x"67800000",
         356 => x"37c50100",
         357 => x"130101f8",
         358 => x"93050000",
         359 => x"13050520",
         360 => x"232e1106",
         361 => x"232c8106",
         362 => x"232a9106",
         363 => x"23282107",
         364 => x"23263107",
         365 => x"23244107",
         366 => x"23225107",
         367 => x"23206107",
         368 => x"232e7105",
         369 => x"232c8105",
         370 => x"232a9105",
         371 => x"2328a105",
         372 => x"2326b105",
         373 => x"eff09fcc",
         374 => x"37150010",
         375 => x"130505c0",
         376 => x"eff09fd0",
         377 => x"37150010",
         378 => x"130545c2",
         379 => x"eff0dfcf",
         380 => x"732510fc",
         381 => x"37190010",
         382 => x"eff0dfe9",
         383 => x"130509c2",
         384 => x"eff09fce",
         385 => x"b70700f0",
         386 => x"1307f03f",
         387 => x"370a1000",
         388 => x"b709a000",
         389 => x"23a2e700",
         390 => x"93041000",
         391 => x"130afaff",
         392 => x"b70a00f0",
         393 => x"93891900",
         394 => x"b3f74401",
         395 => x"639c0700",
         396 => x"1305a002",
         397 => x"eff05fc9",
         398 => x"83a74a00",
         399 => x"93d71700",
         400 => x"23a2fa00",
         401 => x"eff01faa",
         402 => x"13040500",
         403 => x"631a050c",
         404 => x"93841400",
         405 => x"e39a34fd",
         406 => x"b70700f0",
         407 => x"23a20700",
         408 => x"631a0400",
         409 => x"93050000",
         410 => x"13050000",
         411 => x"eff01fc3",
         412 => x"e7000400",
         413 => x"eff01fa8",
         414 => x"93071002",
         415 => x"93040000",
         416 => x"631cf51c",
         417 => x"37140010",
         418 => x"130584c3",
         419 => x"eff0dfc5",
         420 => x"b70900f0",
         421 => x"930a3005",
         422 => x"130ba004",
         423 => x"930b3002",
         424 => x"130a2000",
         425 => x"130ca000",
         426 => x"83a74900",
         427 => x"93c71700",
         428 => x"23a2f900",
         429 => x"eff01fa4",
         430 => x"1375f50f",
         431 => x"63185517",
         432 => x"eff05fa3",
         433 => x"937cf50f",
         434 => x"9387fcfc",
         435 => x"93f7f70f",
         436 => x"6360fa10",
         437 => x"93071003",
         438 => x"6398fc04",
         439 => x"13052000",
         440 => x"eff09fc4",
         441 => x"130dd5ff",
         442 => x"13054000",
         443 => x"eff0dfc3",
         444 => x"b70d01ff",
         445 => x"930c0500",
         446 => x"330dad00",
         447 => x"938dfdff",
         448 => x"639aac05",
         449 => x"930ca000",
         450 => x"eff0df9e",
         451 => x"1375f50f",
         452 => x"e31c95ff",
         453 => x"130584c3",
         454 => x"eff01fbd",
         455 => x"6ff0dff8",
         456 => x"13041000",
         457 => x"6ff05ff3",
         458 => x"93072003",
         459 => x"13052000",
         460 => x"639afc00",
         461 => x"eff05fbf",
         462 => x"130dc5ff",
         463 => x"13056000",
         464 => x"6ff0dffa",
         465 => x"eff05fbe",
         466 => x"130db5ff",
         467 => x"13058000",
         468 => x"6ff0dff9",
         469 => x"93f5ccff",
         470 => x"13052000",
         471 => x"2326b100",
         472 => x"eff09fbc",
         473 => x"8325c100",
         474 => x"93070500",
         475 => x"b7060001",
         476 => x"3706ffff",
         477 => x"13f53c00",
         478 => x"03a70500",
         479 => x"13083000",
         480 => x"9386f6ff",
         481 => x"93081000",
         482 => x"1306f60f",
         483 => x"63064503",
         484 => x"630a0503",
         485 => x"630c1501",
         486 => x"137707f0",
         487 => x"b3e7e700",
         488 => x"23a0f500",
         489 => x"938c1c00",
         490 => x"6ff09ff5",
         491 => x"3377c700",
         492 => x"93978700",
         493 => x"6ff09ffe",
         494 => x"3377b701",
         495 => x"93970701",
         496 => x"6ff0dffd",
         497 => x"3377d700",
         498 => x"93978701",
         499 => x"6ff01ffd",
         500 => x"93879cfc",
         501 => x"93f7f70f",
         502 => x"6362fa04",
         503 => x"13052000",
         504 => x"eff09fb4",
         505 => x"93077003",
         506 => x"13058000",
         507 => x"638afc00",
         508 => x"93078003",
         509 => x"13056000",
         510 => x"6384fc00",
         511 => x"13054000",
         512 => x"eff09fb2",
         513 => x"93040500",
         514 => x"930ca000",
         515 => x"eff09f8e",
         516 => x"1375f50f",
         517 => x"e31c95ff",
         518 => x"6ff0dfef",
         519 => x"eff09f8d",
         520 => x"1375f50f",
         521 => x"e31c85ff",
         522 => x"6ff0dfee",
         523 => x"63186509",
         524 => x"130584c3",
         525 => x"eff05fab",
         526 => x"93050000",
         527 => x"13050000",
         528 => x"eff0dfa5",
         529 => x"23a20900",
         530 => x"e7800400",
         531 => x"b70700f0",
         532 => x"1307a00a",
         533 => x"23a2e700",
         534 => x"130509c2",
         535 => x"b7190010",
         536 => x"eff09fa8",
         537 => x"13040000",
         538 => x"371b0010",
         539 => x"b71b0010",
         540 => x"938959d6",
         541 => x"b7170010",
         542 => x"1385c7c3",
         543 => x"eff0dfa6",
         544 => x"93059002",
         545 => x"13054101",
         546 => x"eff09f88",
         547 => x"13054101",
         548 => x"ef00c02c",
         549 => x"b7170010",
         550 => x"130a0500",
         551 => x"938507c4",
         552 => x"13054101",
         553 => x"eff0df81",
         554 => x"631e0500",
         555 => x"37150010",
         556 => x"130545c4",
         557 => x"eff05fa3",
         558 => x"6f004003",
         559 => x"e31c75e5",
         560 => x"6ff0dff8",
         561 => x"b7170010",
         562 => x"938507d3",
         563 => x"13054101",
         564 => x"eff00fff",
         565 => x"63100502",
         566 => x"93050000",
         567 => x"eff01f9c",
         568 => x"b70700f0",
         569 => x"23a20700",
         570 => x"e7800400",
         571 => x"e3040af8",
         572 => x"6f004018",
         573 => x"b7170010",
         574 => x"13063000",
         575 => x"938547d3",
         576 => x"13054101",
         577 => x"ef004027",
         578 => x"63100504",
         579 => x"93050000",
         580 => x"13057101",
         581 => x"eff09fac",
         582 => x"93773500",
         583 => x"13040500",
         584 => x"63940706",
         585 => x"93058000",
         586 => x"eff0dfbf",
         587 => x"37150010",
         588 => x"130585d3",
         589 => x"eff05f9b",
         590 => x"03250400",
         591 => x"93058000",
         592 => x"eff05fbe",
         593 => x"6ff09ffa",
         594 => x"13063000",
         595 => x"93054bd5",
         596 => x"13054101",
         597 => x"ef004022",
         598 => x"631e0502",
         599 => x"93050101",
         600 => x"13057101",
         601 => x"eff09fa7",
         602 => x"93773500",
         603 => x"13040500",
         604 => x"639c0700",
         605 => x"03250101",
         606 => x"93050000",
         607 => x"eff01fa6",
         608 => x"2320a400",
         609 => x"6ff09ff6",
         610 => x"37150010",
         611 => x"1305c5d3",
         612 => x"6ff05ff2",
         613 => x"13063000",
         614 => x"93858bd5",
         615 => x"13054101",
         616 => x"ef00801d",
         617 => x"83474101",
         618 => x"1307e006",
         619 => x"630c0508",
         620 => x"639ae70a",
         621 => x"93773400",
         622 => x"e39807fc",
         623 => x"130c0404",
         624 => x"b71c0010",
         625 => x"371d0010",
         626 => x"930d80ff",
         627 => x"93058000",
         628 => x"13050400",
         629 => x"eff01fb5",
         630 => x"13858cd3",
         631 => x"eff0df90",
         632 => x"83270400",
         633 => x"93058000",
         634 => x"130a8001",
         635 => x"13850700",
         636 => x"2326f100",
         637 => x"eff01fb3",
         638 => x"1305cdd5",
         639 => x"eff0df8e",
         640 => x"b70a00ff",
         641 => x"8327c100",
         642 => x"33f55701",
         643 => x"33554501",
         644 => x"b3063501",
         645 => x"83c60600",
         646 => x"93f67609",
         647 => x"63800604",
         648 => x"130a8aff",
         649 => x"eff05f8a",
         650 => x"93da8a00",
         651 => x"e31cbafd",
         652 => x"13044400",
         653 => x"130509c2",
         654 => x"eff01f8b",
         655 => x"e31884f9",
         656 => x"6ff05fe3",
         657 => x"e388e7f6",
         658 => x"93050000",
         659 => x"13057101",
         660 => x"eff0df98",
         661 => x"13040500",
         662 => x"6ff0dff5",
         663 => x"1305e002",
         664 => x"6ff01ffc",
         665 => x"e3080ae0",
         666 => x"37150010",
         667 => x"130505d6",
         668 => x"eff09f87",
         669 => x"130509c2",
         670 => x"eff01f87",
         671 => x"6ff09fdf",
         672 => x"130101ff",
         673 => x"23248100",
         674 => x"23261100",
         675 => x"93070000",
         676 => x"13040500",
         677 => x"63880700",
         678 => x"93050000",
         679 => x"97000000",
         680 => x"e7000000",
         681 => x"b7170010",
         682 => x"03a547e7",
         683 => x"83278502",
         684 => x"63840700",
         685 => x"e7800700",
         686 => x"13050400",
         687 => x"eff04fe2",
         688 => x"130101ff",
         689 => x"23248100",
         690 => x"23229100",
         691 => x"37140010",
         692 => x"b7140010",
         693 => x"938784e7",
         694 => x"130484e7",
         695 => x"3304f440",
         696 => x"23202101",
         697 => x"23261100",
         698 => x"13542440",
         699 => x"938484e7",
         700 => x"13090000",
         701 => x"63108904",
         702 => x"b7140010",
         703 => x"37140010",
         704 => x"938784e7",
         705 => x"130484e7",
         706 => x"3304f440",
         707 => x"13542440",
         708 => x"938484e7",
         709 => x"13090000",
         710 => x"63188902",
         711 => x"8320c100",
         712 => x"03248100",
         713 => x"83244100",
         714 => x"03290100",
         715 => x"13010101",
         716 => x"67800000",
         717 => x"83a70400",
         718 => x"13091900",
         719 => x"93844400",
         720 => x"e7800700",
         721 => x"6ff01ffb",
         722 => x"83a70400",
         723 => x"13091900",
         724 => x"93844400",
         725 => x"e7800700",
         726 => x"6ff01ffc",
         727 => x"93070500",
         728 => x"03c70700",
         729 => x"93871700",
         730 => x"e31c07fe",
         731 => x"3385a740",
         732 => x"1305f5ff",
         733 => x"67800000",
         734 => x"630a0602",
         735 => x"1306f6ff",
         736 => x"13070000",
         737 => x"b307e500",
         738 => x"b386e500",
         739 => x"83c70700",
         740 => x"83c60600",
         741 => x"6398d700",
         742 => x"6306c700",
         743 => x"13071700",
         744 => x"e39207fe",
         745 => x"3385d740",
         746 => x"67800000",
         747 => x"13050000",
         748 => x"67800000",
         749 => x"74020010",
         750 => x"b8010010",
         751 => x"b8010010",
         752 => x"b8010010",
         753 => x"b8010010",
         754 => x"18020010",
         755 => x"b8010010",
         756 => x"2c020010",
         757 => x"b8010010",
         758 => x"b8010010",
         759 => x"2c020010",
         760 => x"b8010010",
         761 => x"b8010010",
         762 => x"b8010010",
         763 => x"b8010010",
         764 => x"b8010010",
         765 => x"b8010010",
         766 => x"b8010010",
         767 => x"8c010010",
         768 => x"0d0a5448",
         769 => x"55415320",
         770 => x"52495343",
         771 => x"2d562042",
         772 => x"6f6f746c",
         773 => x"6f616465",
         774 => x"72207630",
         775 => x"2e342e31",
         776 => x"0d0a0000",
         777 => x"436c6f63",
         778 => x"6b206672",
         779 => x"65717565",
         780 => x"6e63793a",
         781 => x"20000000",
         782 => x"3f0a0000",
         783 => x"3e200000",
         784 => x"68000000",
         785 => x"48656c70",
         786 => x"3a0d0a20",
         787 => x"68202020",
         788 => x"20202020",
         789 => x"20202020",
         790 => x"20202020",
         791 => x"202d2074",
         792 => x"68697320",
         793 => x"68656c70",
         794 => x"0d0a2072",
         795 => x"20202020",
         796 => x"20202020",
         797 => x"20202020",
         798 => x"20202020",
         799 => x"2d207275",
         800 => x"6e206170",
         801 => x"706c6963",
         802 => x"6174696f",
         803 => x"6e0d0a20",
         804 => x"7277203c",
         805 => x"61646472",
         806 => x"3e202020",
         807 => x"20202020",
         808 => x"202d2072",
         809 => x"65616420",
         810 => x"776f7264",
         811 => x"2066726f",
         812 => x"6d206164",
         813 => x"64720d0a",
         814 => x"20777720",
         815 => x"3c616464",
         816 => x"723e203c",
         817 => x"64617461",
         818 => x"3e202d20",
         819 => x"77726974",
         820 => x"6520776f",
         821 => x"72642064",
         822 => x"61746120",
         823 => x"61742061",
         824 => x"6464720d",
         825 => x"0a206477",
         826 => x"203c6164",
         827 => x"64723e20",
         828 => x"20202020",
         829 => x"2020202d",
         830 => x"2064756d",
         831 => x"70203136",
         832 => x"20776f72",
         833 => x"64730d0a",
         834 => x"206e2020",
         835 => x"20202020",
         836 => x"20202020",
         837 => x"20202020",
         838 => x"20202d20",
         839 => x"64756d70",
         840 => x"206e6578",
         841 => x"74203136",
         842 => x"20776f72",
         843 => x"64730000",
         844 => x"72000000",
         845 => x"72772000",
         846 => x"3a200000",
         847 => x"4e6f7420",
         848 => x"6f6e2034",
         849 => x"2d627974",
         850 => x"6520626f",
         851 => x"756e6461",
         852 => x"72792100",
         853 => x"77772000",
         854 => x"64772000",
         855 => x"20200000",
         856 => x"3f3f0000",
         857 => x"00202020",
         858 => x"20202020",
         859 => x"20202828",
         860 => x"28282820",
         861 => x"20202020",
         862 => x"20202020",
         863 => x"20202020",
         864 => x"20202020",
         865 => x"20881010",
         866 => x"10101010",
         867 => x"10101010",
         868 => x"10101010",
         869 => x"10040404",
         870 => x"04040404",
         871 => x"04040410",
         872 => x"10101010",
         873 => x"10104141",
         874 => x"41414141",
         875 => x"01010101",
         876 => x"01010101",
         877 => x"01010101",
         878 => x"01010101",
         879 => x"01010101",
         880 => x"10101010",
         881 => x"10104242",
         882 => x"42424242",
         883 => x"02020202",
         884 => x"02020202",
         885 => x"02020202",
         886 => x"02020202",
         887 => x"02020202",
         888 => x"10101010",
         889 => x"20000000",
         890 => x"00000000",
         891 => x"00000000",
         892 => x"00000000",
         893 => x"00000000",
         894 => x"00000000",
         895 => x"00000000",
         896 => x"00000000",
         897 => x"00000000",
         898 => x"00000000",
         899 => x"00000000",
         900 => x"00000000",
         901 => x"00000000",
         902 => x"00000000",
         903 => x"00000000",
         904 => x"00000000",
         905 => x"00000000",
         906 => x"00000000",
         907 => x"00000000",
         908 => x"00000000",
         909 => x"00000000",
         910 => x"00000000",
         911 => x"00000000",
         912 => x"00000000",
         913 => x"00000000",
         914 => x"00000000",
         915 => x"00000000",
         916 => x"00000000",
         917 => x"00000000",
         918 => x"00000000",
         919 => x"00000000",
         920 => x"00000000",
         921 => x"00000000",
         922 => x"3c627265",
         923 => x"616b3e0d",
         924 => x"0a000000",
         925 => x"00000020",
         926 => x"00000000",
         927 => x"00000000",
         928 => x"00000000",
         929 => x"00000000",
         930 => x"00000000",
         931 => x"00000000",
         932 => x"00000000",
         933 => x"00000000",
         934 => x"00000000",
         935 => x"00000000",
         936 => x"00000000",
         937 => x"00000000",
         938 => x"00000000",
         939 => x"00000000",
         940 => x"00000000",
         941 => x"00000000",
         942 => x"00000000",
         943 => x"00000000",
         944 => x"00000000",
         945 => x"00000000",
         946 => x"00000000",
         947 => x"00000000",
         948 => x"00000000",
         949 => x"00000000",
         950 => x"00000020",
         others => (others => '0')
        );

begin

    gen_bootrom: if HAVE_BOOTLOADER_ROM generate

        -- ROM, for both instructions and read-only data
        process (I_clk, I_areset, I_pc, I_memaddress, I_csboot, I_memsize, I_stall) is
        variable address_instr : integer range 0 to bootloader_size-1;
        variable address_data : integer range 0 to bootloader_size-1;
        variable instr_var : data_type;
        variable instr_recode : data_type;
        variable romdata_var : data_type;
        constant x : data_type := (others => 'X');
        begin
            -- Calculate addresses
            address_instr := to_integer(unsigned(I_pc(bootloader_size_bits-1 downto 2)));
            address_data := to_integer(unsigned(I_memaddress(bootloader_size_bits-1 downto 2)));

            -- Quartus will detect ROM table and uses onboard RAM
            -- Do not use reset, otherwise ROM will be created with ALMs
            if rising_edge(I_clk) then
                if I_stall = '0' then
                    instr_var := bootrom(address_instr);
                end if;
                romdata_var := bootrom(address_data);
            end if;
            
            -- Recode instruction
            O_instr <= instr_var(7 downto 0) & instr_var(15 downto 8) & instr_var(23 downto 16) & instr_var(31 downto 24);
            
            O_load_misaligned_error <= '0';
            
            -- By natural size, for data
            if I_csboot = '1' then
                if I_memsize = memsize_word and I_memaddress(1 downto 0) = "00" then
                    O_dataout <= romdata_var(7 downto 0) & romdata_var(15 downto 8) & romdata_var(23 downto 16) & romdata_var(31 downto 24);
                elsif I_memsize = memsize_halfword and I_memaddress(1 downto 0) = "00" then
                    O_dataout <= x(31 downto 16) & romdata_var(23 downto 16) & romdata_var(31 downto 24);
                elsif I_memsize = memsize_halfword and I_memaddress(1 downto 0) = "10" then
                    O_dataout <= x(31 downto 16) & romdata_var(7 downto 0) & romdata_var(15 downto 8);
                elsif I_memsize = memsize_byte then
                    case I_memaddress(1 downto 0) is
                        when "00" => O_dataout <= x(31 downto 8) & romdata_var(31 downto 24);
                        when "01" => O_dataout <= x(31 downto 8) & romdata_var(23 downto 16);
                        when "10" => O_dataout <= x(31 downto 8) & romdata_var(15 downto 8);
                        when "11" => O_dataout <= x(31 downto 8) & romdata_var(7 downto 0);
                        when others => O_dataout <= x; O_load_misaligned_error <= '1';
                    end case;
                else
                    -- Chip select, but not aligned
                    O_dataout <= x;
                    O_load_misaligned_error <= '1';
                end if;
            else
                -- No chip select, so no data
                O_dataout <= x;
            end if;
        end process;
    end generate;

    gen_bootrom_not: if not HAVE_BOOTLOADER_ROM generate
        O_load_misaligned_error <= '0';
        O_dataout <= (others => 'X');
        O_instr  <= (others => 'X');
    end generate;
end architecture rtl;
