-- srec2vhdl table generator
-- for input file 'interrupt_direct.srec'
-- date: Sun May 21 14:32:29 2023


library ieee;
use ieee.std_logic_1164.all;

library work;
use work.processor_common.all;

package processor_common_rom is
    constant rom_contents : rom_type := (
           0 => x"97020000",
           1 => x"93820228",
           2 => x"73905230",
           3 => x"97010020",
           4 => x"9381417f",
           5 => x"17810020",
           6 => x"1301c1fe",
           7 => x"13860188",
           8 => x"93874189",
           9 => x"637af600",
          10 => x"3386c740",
          11 => x"93050000",
          12 => x"13850188",
          13 => x"ef108030",
          14 => x"37050020",
          15 => x"13060500",
          16 => x"93870188",
          17 => x"637cf600",
          18 => x"b7350000",
          19 => x"3386c740",
          20 => x"9385c502",
          21 => x"13050500",
          22 => x"ef10002c",
          23 => x"ef10d002",
          24 => x"b7050020",
          25 => x"13060000",
          26 => x"93850500",
          27 => x"13055000",
          28 => x"ef10404c",
          29 => x"ef10407d",
          30 => x"6f104041",
          31 => x"130101ff",
          32 => x"23261100",
          33 => x"ef100045",
          34 => x"8320c100",
          35 => x"13051000",
          36 => x"13010101",
          37 => x"67800000",
          38 => x"130101fd",
          39 => x"232c4101",
          40 => x"130a0500",
          41 => x"37350000",
          42 => x"130585e7",
          43 => x"23248102",
          44 => x"23229102",
          45 => x"23202103",
          46 => x"232e3101",
          47 => x"83244a08",
          48 => x"23261102",
          49 => x"13044100",
          50 => x"ef10c042",
          51 => x"37390000",
          52 => x"9309c1ff",
          53 => x"93070400",
          54 => x"1309c9c4",
          55 => x"13f7f400",
          56 => x"3307e900",
          57 => x"03470700",
          58 => x"9387f7ff",
          59 => x"93d44400",
          60 => x"2384e700",
          61 => x"e39437ff",
          62 => x"13054100",
          63 => x"23060100",
          64 => x"ef10403f",
          65 => x"37350000",
          66 => x"1305c5e8",
          67 => x"ef10803e",
          68 => x"03278a08",
          69 => x"9377f700",
          70 => x"b307f900",
          71 => x"83c70700",
          72 => x"1304f4ff",
          73 => x"13574700",
          74 => x"2304f400",
          75 => x"e31434ff",
          76 => x"13054100",
          77 => x"ef10003c",
          78 => x"37350000",
          79 => x"130545ec",
          80 => x"ef10403b",
          81 => x"8320c102",
          82 => x"03248102",
          83 => x"83244102",
          84 => x"03290102",
          85 => x"8329c101",
          86 => x"032a8101",
          87 => x"13010103",
          88 => x"67800000",
          89 => x"b70700f0",
          90 => x"03a74708",
          91 => x"1377f7fe",
          92 => x"23a2e708",
          93 => x"03a74700",
          94 => x"13471700",
          95 => x"23a2e700",
          96 => x"67800000",
          97 => x"370700f0",
          98 => x"83274700",
          99 => x"93e70720",
         100 => x"2322f700",
         101 => x"6f000000",
         102 => x"b70700f0",
         103 => x"83a6470f",
         104 => x"03a6070f",
         105 => x"03a7470f",
         106 => x"e31ad7fe",
         107 => x"b7860100",
         108 => x"9305f0ff",
         109 => x"9386066a",
         110 => x"23aeb70e",
         111 => x"b306d600",
         112 => x"23acb70e",
         113 => x"33b6c600",
         114 => x"23acd70e",
         115 => x"3306e600",
         116 => x"23aec70e",
         117 => x"03a74700",
         118 => x"13472700",
         119 => x"23a2e700",
         120 => x"67800000",
         121 => x"b70700f0",
         122 => x"03a74702",
         123 => x"13774700",
         124 => x"630a0700",
         125 => x"03a74700",
         126 => x"13478700",
         127 => x"23a2e700",
         128 => x"83a78702",
         129 => x"67800000",
         130 => x"b70700f0",
         131 => x"03a7470a",
         132 => x"1377f7f0",
         133 => x"23a2e70a",
         134 => x"03a74700",
         135 => x"13474700",
         136 => x"23a2e700",
         137 => x"67800000",
         138 => x"b70700f0",
         139 => x"03a74706",
         140 => x"137777ff",
         141 => x"23a2e706",
         142 => x"03a74700",
         143 => x"13470701",
         144 => x"23a2e700",
         145 => x"67800000",
         146 => x"b70700f0",
         147 => x"03a74704",
         148 => x"137777fe",
         149 => x"23a2e704",
         150 => x"03a74700",
         151 => x"13470702",
         152 => x"23a2e700",
         153 => x"67800000",
         154 => x"b70700f0",
         155 => x"23ae0700",
         156 => x"03a74700",
         157 => x"13470704",
         158 => x"23a2e700",
         159 => x"67800000",
         160 => x"6f000000",
         161 => x"13050000",
         162 => x"67800000",
         163 => x"13050000",
         164 => x"67800000",
         165 => x"130101f7",
         166 => x"23221100",
         167 => x"23242100",
         168 => x"23263100",
         169 => x"23284100",
         170 => x"232a5100",
         171 => x"232c6100",
         172 => x"232e7100",
         173 => x"23208102",
         174 => x"23229102",
         175 => x"2324a102",
         176 => x"2326b102",
         177 => x"2328c102",
         178 => x"232ad102",
         179 => x"232ce102",
         180 => x"232ef102",
         181 => x"23200105",
         182 => x"23221105",
         183 => x"23242105",
         184 => x"23263105",
         185 => x"23284105",
         186 => x"232a5105",
         187 => x"232c6105",
         188 => x"232e7105",
         189 => x"23208107",
         190 => x"23229107",
         191 => x"2324a107",
         192 => x"2326b107",
         193 => x"2328c107",
         194 => x"232ad107",
         195 => x"232ce107",
         196 => x"232ef107",
         197 => x"f3222034",
         198 => x"23205108",
         199 => x"f3221034",
         200 => x"23225108",
         201 => x"83a20200",
         202 => x"23245108",
         203 => x"f3223034",
         204 => x"23265108",
         205 => x"f3272034",
         206 => x"37070080",
         207 => x"93067700",
         208 => x"6380d710",
         209 => x"9306b000",
         210 => x"63fef602",
         211 => x"934607ff",
         212 => x"b386d700",
         213 => x"13065000",
         214 => x"636ad602",
         215 => x"1347f7fe",
         216 => x"b387e700",
         217 => x"13074000",
         218 => x"6364f716",
         219 => x"37370000",
         220 => x"93972700",
         221 => x"130707c6",
         222 => x"b387e700",
         223 => x"83a70700",
         224 => x"67800700",
         225 => x"13071000",
         226 => x"636ef708",
         227 => x"03258102",
         228 => x"83220108",
         229 => x"63c80200",
         230 => x"f3221034",
         231 => x"93824200",
         232 => x"73901234",
         233 => x"832fc107",
         234 => x"032f8107",
         235 => x"832e4107",
         236 => x"032e0107",
         237 => x"832dc106",
         238 => x"032d8106",
         239 => x"832c4106",
         240 => x"032c0106",
         241 => x"832bc105",
         242 => x"032b8105",
         243 => x"832a4105",
         244 => x"032a0105",
         245 => x"8329c104",
         246 => x"03298104",
         247 => x"83284104",
         248 => x"03280104",
         249 => x"8327c103",
         250 => x"03278103",
         251 => x"83264103",
         252 => x"03260103",
         253 => x"8325c102",
         254 => x"83244102",
         255 => x"03240102",
         256 => x"8323c101",
         257 => x"03238101",
         258 => x"83224101",
         259 => x"03220101",
         260 => x"8321c100",
         261 => x"03218100",
         262 => x"83204100",
         263 => x"13010109",
         264 => x"73002030",
         265 => x"e3e4f6f6",
         266 => x"37370000",
         267 => x"93972700",
         268 => x"130747c7",
         269 => x"b387e700",
         270 => x"83a70700",
         271 => x"67800700",
         272 => x"eff09fd5",
         273 => x"03258102",
         274 => x"6ff09ff4",
         275 => x"eff0dfdb",
         276 => x"03258102",
         277 => x"6ff0dff3",
         278 => x"eff01fdd",
         279 => x"03258102",
         280 => x"6ff01ff3",
         281 => x"eff05fde",
         282 => x"03258102",
         283 => x"6ff05ff2",
         284 => x"eff05fcf",
         285 => x"03258102",
         286 => x"6ff09ff1",
         287 => x"eff09fd6",
         288 => x"03258102",
         289 => x"6ff0dff0",
         290 => x"9307600d",
         291 => x"6384f806",
         292 => x"9307900a",
         293 => x"6388f818",
         294 => x"63ca170f",
         295 => x"938878fc",
         296 => x"93074002",
         297 => x"63ec1703",
         298 => x"b7370000",
         299 => x"938747ca",
         300 => x"93982800",
         301 => x"b388f800",
         302 => x"83a70800",
         303 => x"67800700",
         304 => x"13050100",
         305 => x"eff05fbd",
         306 => x"03258102",
         307 => x"6ff05fec",
         308 => x"eff09fd9",
         309 => x"03258102",
         310 => x"6ff09feb",
         311 => x"ef104036",
         312 => x"93078005",
         313 => x"2320f500",
         314 => x"9307f0ff",
         315 => x"13850700",
         316 => x"6ff01fea",
         317 => x"63120510",
         318 => x"13858189",
         319 => x"13050500",
         320 => x"6ff01fe9",
         321 => x"b7270000",
         322 => x"23a2f500",
         323 => x"93070000",
         324 => x"13850700",
         325 => x"6ff0dfe7",
         326 => x"93070000",
         327 => x"13850700",
         328 => x"6ff01fe7",
         329 => x"ef10c031",
         330 => x"93079000",
         331 => x"2320f500",
         332 => x"9307f0ff",
         333 => x"13850700",
         334 => x"6ff09fe5",
         335 => x"13090600",
         336 => x"13840500",
         337 => x"635cc000",
         338 => x"b384c500",
         339 => x"03450400",
         340 => x"13041400",
         341 => x"eff09fb2",
         342 => x"e39a84fe",
         343 => x"13050900",
         344 => x"6ff01fe3",
         345 => x"13090600",
         346 => x"13840500",
         347 => x"e358c0fe",
         348 => x"b384c500",
         349 => x"eff05fb0",
         350 => x"2300a400",
         351 => x"13041400",
         352 => x"e31a94fe",
         353 => x"13050900",
         354 => x"6ff09fe0",
         355 => x"938808c0",
         356 => x"9307f000",
         357 => x"e3e417f5",
         358 => x"b7370000",
         359 => x"938787d3",
         360 => x"93982800",
         361 => x"b388f800",
         362 => x"83a70800",
         363 => x"67800700",
         364 => x"ef100029",
         365 => x"9307d000",
         366 => x"2320f500",
         367 => x"9307f0ff",
         368 => x"13850700",
         369 => x"6ff0dfdc",
         370 => x"ef108027",
         371 => x"93072000",
         372 => x"2320f500",
         373 => x"9307f0ff",
         374 => x"13850700",
         375 => x"6ff05fdb",
         376 => x"ef100026",
         377 => x"9307f001",
         378 => x"2320f500",
         379 => x"9307f0ff",
         380 => x"13850700",
         381 => x"6ff0dfd9",
         382 => x"b7870020",
         383 => x"93870700",
         384 => x"13070040",
         385 => x"b387e740",
         386 => x"e36af5ee",
         387 => x"ef104023",
         388 => x"9307c000",
         389 => x"2320f500",
         390 => x"1305f0ff",
         391 => x"13050500",
         392 => x"6ff01fd7",
         393 => x"13090000",
         394 => x"93040500",
         395 => x"13040900",
         396 => x"93090900",
         397 => x"93070900",
         398 => x"732410c8",
         399 => x"f32910c0",
         400 => x"f32710c8",
         401 => x"e31af4fe",
         402 => x"37460f00",
         403 => x"13060624",
         404 => x"93060000",
         405 => x"13850900",
         406 => x"93050400",
         407 => x"ef00900d",
         408 => x"37460f00",
         409 => x"23a4a400",
         410 => x"13060624",
         411 => x"93060000",
         412 => x"13850900",
         413 => x"93050400",
         414 => x"ef00c048",
         415 => x"23a0a400",
         416 => x"23a2b400",
         417 => x"13050900",
         418 => x"6ff09fd0",
         419 => x"13030500",
         420 => x"138e0500",
         421 => x"93080000",
         422 => x"63dc0500",
         423 => x"b337a000",
         424 => x"330eb040",
         425 => x"330efe40",
         426 => x"3303a040",
         427 => x"9308f0ff",
         428 => x"63dc0600",
         429 => x"b337c000",
         430 => x"b306d040",
         431 => x"93c8f8ff",
         432 => x"b386f640",
         433 => x"3306c040",
         434 => x"13070600",
         435 => x"13080300",
         436 => x"93070e00",
         437 => x"639c0628",
         438 => x"b7350000",
         439 => x"938585d7",
         440 => x"6376ce0e",
         441 => x"b7060100",
         442 => x"6378d60c",
         443 => x"93360610",
         444 => x"93c61600",
         445 => x"93963600",
         446 => x"3355d600",
         447 => x"b385a500",
         448 => x"83c50500",
         449 => x"13050002",
         450 => x"b386d500",
         451 => x"b305d540",
         452 => x"630cd500",
         453 => x"b317be00",
         454 => x"b356d300",
         455 => x"3317b600",
         456 => x"b3e7f600",
         457 => x"3318b300",
         458 => x"93550701",
         459 => x"33deb702",
         460 => x"13160701",
         461 => x"13560601",
         462 => x"b3f7b702",
         463 => x"13050e00",
         464 => x"3303c603",
         465 => x"93960701",
         466 => x"93570801",
         467 => x"b3e7d700",
         468 => x"63fe6700",
         469 => x"b307f700",
         470 => x"1305feff",
         471 => x"63e8e700",
         472 => x"63f66700",
         473 => x"1305eeff",
         474 => x"b387e700",
         475 => x"b3876740",
         476 => x"33d3b702",
         477 => x"13180801",
         478 => x"13580801",
         479 => x"b3f7b702",
         480 => x"b3066602",
         481 => x"93970701",
         482 => x"3368f800",
         483 => x"93070300",
         484 => x"637cd800",
         485 => x"33080701",
         486 => x"9307f3ff",
         487 => x"6366e800",
         488 => x"6374d800",
         489 => x"9307e3ff",
         490 => x"13150501",
         491 => x"3365f500",
         492 => x"93050000",
         493 => x"6f00000e",
         494 => x"37050001",
         495 => x"93060001",
         496 => x"e36ca6f2",
         497 => x"93068001",
         498 => x"6ff01ff3",
         499 => x"93060000",
         500 => x"630c0600",
         501 => x"b7070100",
         502 => x"637af60c",
         503 => x"93360610",
         504 => x"93c61600",
         505 => x"93963600",
         506 => x"b357d600",
         507 => x"b385f500",
         508 => x"83c70500",
         509 => x"b387d700",
         510 => x"93060002",
         511 => x"b385f640",
         512 => x"6390f60c",
         513 => x"b307ce40",
         514 => x"93051000",
         515 => x"13530701",
         516 => x"b3de6702",
         517 => x"13160701",
         518 => x"13560601",
         519 => x"93560801",
         520 => x"b3f76702",
         521 => x"13850e00",
         522 => x"330ed603",
         523 => x"93970701",
         524 => x"b3e7f600",
         525 => x"63fec701",
         526 => x"b307f700",
         527 => x"1385feff",
         528 => x"63e8e700",
         529 => x"63f6c701",
         530 => x"1385eeff",
         531 => x"b387e700",
         532 => x"b387c741",
         533 => x"33de6702",
         534 => x"13180801",
         535 => x"13580801",
         536 => x"b3f76702",
         537 => x"b306c603",
         538 => x"93970701",
         539 => x"3368f800",
         540 => x"93070e00",
         541 => x"637cd800",
         542 => x"33080701",
         543 => x"9307feff",
         544 => x"6366e800",
         545 => x"6374d800",
         546 => x"9307eeff",
         547 => x"13150501",
         548 => x"3365f500",
         549 => x"638a0800",
         550 => x"b337a000",
         551 => x"b305b040",
         552 => x"b385f540",
         553 => x"3305a040",
         554 => x"67800000",
         555 => x"b7070001",
         556 => x"93060001",
         557 => x"e36af6f2",
         558 => x"93068001",
         559 => x"6ff0dff2",
         560 => x"3317b600",
         561 => x"b356fe00",
         562 => x"13550701",
         563 => x"331ebe00",
         564 => x"b357f300",
         565 => x"b3e7c701",
         566 => x"33dea602",
         567 => x"13160701",
         568 => x"13560601",
         569 => x"3318b300",
         570 => x"b3f6a602",
         571 => x"3303c603",
         572 => x"93950601",
         573 => x"93d60701",
         574 => x"b3e6b600",
         575 => x"93050e00",
         576 => x"63fe6600",
         577 => x"b306d700",
         578 => x"9305feff",
         579 => x"63e8e600",
         580 => x"63f66600",
         581 => x"9305eeff",
         582 => x"b386e600",
         583 => x"b3866640",
         584 => x"33d3a602",
         585 => x"93970701",
         586 => x"93d70701",
         587 => x"b3f6a602",
         588 => x"33066602",
         589 => x"93960601",
         590 => x"b3e7d700",
         591 => x"93060300",
         592 => x"63fec700",
         593 => x"b307f700",
         594 => x"9306f3ff",
         595 => x"63e8e700",
         596 => x"63f6c700",
         597 => x"9306e3ff",
         598 => x"b387e700",
         599 => x"93950501",
         600 => x"b387c740",
         601 => x"b3e5d500",
         602 => x"6ff05fea",
         603 => x"6366de18",
         604 => x"b7070100",
         605 => x"63f4f604",
         606 => x"13b70610",
         607 => x"13471700",
         608 => x"13173700",
         609 => x"b7370000",
         610 => x"b3d5e600",
         611 => x"938787d7",
         612 => x"b387b700",
         613 => x"83c70700",
         614 => x"b387e700",
         615 => x"13070002",
         616 => x"b305f740",
         617 => x"6316f702",
         618 => x"13051000",
         619 => x"e3e4c6ef",
         620 => x"3335c300",
         621 => x"13451500",
         622 => x"6ff0dfed",
         623 => x"b7070001",
         624 => x"13070001",
         625 => x"e3e0f6fc",
         626 => x"13078001",
         627 => x"6ff09ffb",
         628 => x"3357f600",
         629 => x"b396b600",
         630 => x"b366d700",
         631 => x"3357fe00",
         632 => x"331ebe00",
         633 => x"b357f300",
         634 => x"b3e7c701",
         635 => x"13de0601",
         636 => x"335fc703",
         637 => x"13980601",
         638 => x"13580801",
         639 => x"3316b600",
         640 => x"3377c703",
         641 => x"b30ee803",
         642 => x"13150701",
         643 => x"13d70701",
         644 => x"3367a700",
         645 => x"13050f00",
         646 => x"637ed701",
         647 => x"3387e600",
         648 => x"1305ffff",
         649 => x"6368d700",
         650 => x"6376d701",
         651 => x"1305efff",
         652 => x"3307d700",
         653 => x"3307d741",
         654 => x"b35ec703",
         655 => x"93970701",
         656 => x"93d70701",
         657 => x"3377c703",
         658 => x"3308d803",
         659 => x"13170701",
         660 => x"b3e7e700",
         661 => x"13870e00",
         662 => x"63fe0701",
         663 => x"b387f600",
         664 => x"1387feff",
         665 => x"63e8d700",
         666 => x"63f60701",
         667 => x"1387eeff",
         668 => x"b387d700",
         669 => x"13150501",
         670 => x"b70e0100",
         671 => x"3365e500",
         672 => x"9386feff",
         673 => x"3377d500",
         674 => x"b3870741",
         675 => x"b376d600",
         676 => x"13580501",
         677 => x"13560601",
         678 => x"330ed702",
         679 => x"b306d802",
         680 => x"3307c702",
         681 => x"3308c802",
         682 => x"3306d700",
         683 => x"13570e01",
         684 => x"3307c700",
         685 => x"6374d700",
         686 => x"3308d801",
         687 => x"93560701",
         688 => x"b3860601",
         689 => x"63e6d702",
         690 => x"e394d7ce",
         691 => x"b7070100",
         692 => x"9387f7ff",
         693 => x"3377f700",
         694 => x"13170701",
         695 => x"337efe00",
         696 => x"3313b300",
         697 => x"3307c701",
         698 => x"93050000",
         699 => x"e374e3da",
         700 => x"1305f5ff",
         701 => x"6ff0dfcb",
         702 => x"93050000",
         703 => x"13050000",
         704 => x"6ff05fd9",
         705 => x"93080500",
         706 => x"13830500",
         707 => x"13070600",
         708 => x"13080500",
         709 => x"93870500",
         710 => x"63920628",
         711 => x"b7350000",
         712 => x"938585d7",
         713 => x"6376c30e",
         714 => x"b7060100",
         715 => x"6378d60c",
         716 => x"93360610",
         717 => x"93c61600",
         718 => x"93963600",
         719 => x"3355d600",
         720 => x"b385a500",
         721 => x"83c50500",
         722 => x"13050002",
         723 => x"b386d500",
         724 => x"b305d540",
         725 => x"630cd500",
         726 => x"b317b300",
         727 => x"b3d6d800",
         728 => x"3317b600",
         729 => x"b3e7f600",
         730 => x"3398b800",
         731 => x"93550701",
         732 => x"33d3b702",
         733 => x"13160701",
         734 => x"13560601",
         735 => x"b3f7b702",
         736 => x"13050300",
         737 => x"b3086602",
         738 => x"93960701",
         739 => x"93570801",
         740 => x"b3e7d700",
         741 => x"63fe1701",
         742 => x"b307f700",
         743 => x"1305f3ff",
         744 => x"63e8e700",
         745 => x"63f61701",
         746 => x"1305e3ff",
         747 => x"b387e700",
         748 => x"b3871741",
         749 => x"b3d8b702",
         750 => x"13180801",
         751 => x"13580801",
         752 => x"b3f7b702",
         753 => x"b3061603",
         754 => x"93970701",
         755 => x"3368f800",
         756 => x"93870800",
         757 => x"637cd800",
         758 => x"33080701",
         759 => x"9387f8ff",
         760 => x"6366e800",
         761 => x"6374d800",
         762 => x"9387e8ff",
         763 => x"13150501",
         764 => x"3365f500",
         765 => x"93050000",
         766 => x"67800000",
         767 => x"37050001",
         768 => x"93060001",
         769 => x"e36ca6f2",
         770 => x"93068001",
         771 => x"6ff01ff3",
         772 => x"93060000",
         773 => x"630c0600",
         774 => x"b7070100",
         775 => x"6370f60c",
         776 => x"93360610",
         777 => x"93c61600",
         778 => x"93963600",
         779 => x"b357d600",
         780 => x"b385f500",
         781 => x"83c70500",
         782 => x"b387d700",
         783 => x"93060002",
         784 => x"b385f640",
         785 => x"6396f60a",
         786 => x"b307c340",
         787 => x"93051000",
         788 => x"93580701",
         789 => x"33de1703",
         790 => x"13160701",
         791 => x"13560601",
         792 => x"93560801",
         793 => x"b3f71703",
         794 => x"13050e00",
         795 => x"3303c603",
         796 => x"93970701",
         797 => x"b3e7f600",
         798 => x"63fe6700",
         799 => x"b307f700",
         800 => x"1305feff",
         801 => x"63e8e700",
         802 => x"63f66700",
         803 => x"1305eeff",
         804 => x"b387e700",
         805 => x"b3876740",
         806 => x"33d31703",
         807 => x"13180801",
         808 => x"13580801",
         809 => x"b3f71703",
         810 => x"b3066602",
         811 => x"93970701",
         812 => x"3368f800",
         813 => x"93070300",
         814 => x"637cd800",
         815 => x"33080701",
         816 => x"9307f3ff",
         817 => x"6366e800",
         818 => x"6374d800",
         819 => x"9307e3ff",
         820 => x"13150501",
         821 => x"3365f500",
         822 => x"67800000",
         823 => x"b7070001",
         824 => x"93060001",
         825 => x"e364f6f4",
         826 => x"93068001",
         827 => x"6ff01ff4",
         828 => x"3317b600",
         829 => x"b356f300",
         830 => x"13550701",
         831 => x"3313b300",
         832 => x"b3d7f800",
         833 => x"b3e76700",
         834 => x"33d3a602",
         835 => x"13160701",
         836 => x"13560601",
         837 => x"3398b800",
         838 => x"b3f6a602",
         839 => x"b3086602",
         840 => x"93950601",
         841 => x"93d60701",
         842 => x"b3e6b600",
         843 => x"93050300",
         844 => x"63fe1601",
         845 => x"b306d700",
         846 => x"9305f3ff",
         847 => x"63e8e600",
         848 => x"63f61601",
         849 => x"9305e3ff",
         850 => x"b386e600",
         851 => x"b3861641",
         852 => x"b3d8a602",
         853 => x"93970701",
         854 => x"93d70701",
         855 => x"b3f6a602",
         856 => x"33061603",
         857 => x"93960601",
         858 => x"b3e7d700",
         859 => x"93860800",
         860 => x"63fec700",
         861 => x"b307f700",
         862 => x"9386f8ff",
         863 => x"63e8e700",
         864 => x"63f6c700",
         865 => x"9386e8ff",
         866 => x"b387e700",
         867 => x"93950501",
         868 => x"b387c740",
         869 => x"b3e5d500",
         870 => x"6ff09feb",
         871 => x"63e6d518",
         872 => x"b7070100",
         873 => x"63f4f604",
         874 => x"13b70610",
         875 => x"13471700",
         876 => x"13173700",
         877 => x"b7370000",
         878 => x"b3d5e600",
         879 => x"938787d7",
         880 => x"b387b700",
         881 => x"83c70700",
         882 => x"b387e700",
         883 => x"13070002",
         884 => x"b305f740",
         885 => x"6316f702",
         886 => x"13051000",
         887 => x"e3ee66e0",
         888 => x"33b5c800",
         889 => x"13451500",
         890 => x"67800000",
         891 => x"b7070001",
         892 => x"13070001",
         893 => x"e3e0f6fc",
         894 => x"13078001",
         895 => x"6ff09ffb",
         896 => x"3357f600",
         897 => x"b396b600",
         898 => x"b366d700",
         899 => x"3357f300",
         900 => x"3313b300",
         901 => x"b3d7f800",
         902 => x"b3e76700",
         903 => x"13d30601",
         904 => x"b35e6702",
         905 => x"13980601",
         906 => x"13580801",
         907 => x"3316b600",
         908 => x"33776702",
         909 => x"330ed803",
         910 => x"13150701",
         911 => x"13d70701",
         912 => x"3367a700",
         913 => x"13850e00",
         914 => x"637ec701",
         915 => x"3387e600",
         916 => x"1385feff",
         917 => x"6368d700",
         918 => x"6376c701",
         919 => x"1385eeff",
         920 => x"3307d700",
         921 => x"3307c741",
         922 => x"335e6702",
         923 => x"93970701",
         924 => x"93d70701",
         925 => x"33776702",
         926 => x"3308c803",
         927 => x"13170701",
         928 => x"b3e7e700",
         929 => x"13070e00",
         930 => x"63fe0701",
         931 => x"b387f600",
         932 => x"1307feff",
         933 => x"63e8d700",
         934 => x"63f60701",
         935 => x"1307eeff",
         936 => x"b387d700",
         937 => x"13150501",
         938 => x"370e0100",
         939 => x"3365e500",
         940 => x"9306feff",
         941 => x"3377d500",
         942 => x"b3870741",
         943 => x"b376d600",
         944 => x"13580501",
         945 => x"13560601",
         946 => x"3303d702",
         947 => x"b306d802",
         948 => x"3307c702",
         949 => x"3308c802",
         950 => x"3306d700",
         951 => x"13570301",
         952 => x"3307c700",
         953 => x"6374d700",
         954 => x"3308c801",
         955 => x"93560701",
         956 => x"b3860601",
         957 => x"63e6d702",
         958 => x"e39ed7ce",
         959 => x"b7070100",
         960 => x"9387f7ff",
         961 => x"3377f700",
         962 => x"13170701",
         963 => x"3373f300",
         964 => x"b398b800",
         965 => x"33076700",
         966 => x"93050000",
         967 => x"e3fee8cc",
         968 => x"1305f5ff",
         969 => x"6ff01fcd",
         970 => x"93050000",
         971 => x"13050000",
         972 => x"67800000",
         973 => x"13080600",
         974 => x"93070500",
         975 => x"13870500",
         976 => x"63960620",
         977 => x"b7380000",
         978 => x"938888d7",
         979 => x"63fcc50c",
         980 => x"b7060100",
         981 => x"637ed60a",
         982 => x"93360610",
         983 => x"93c61600",
         984 => x"93963600",
         985 => x"3353d600",
         986 => x"b3886800",
         987 => x"83c80800",
         988 => x"13030002",
         989 => x"b386d800",
         990 => x"b308d340",
         991 => x"630cd300",
         992 => x"33971501",
         993 => x"b356d500",
         994 => x"33181601",
         995 => x"33e7e600",
         996 => x"b3171501",
         997 => x"13560801",
         998 => x"b356c702",
         999 => x"13150801",
        1000 => x"13550501",
        1001 => x"3377c702",
        1002 => x"b386a602",
        1003 => x"93150701",
        1004 => x"13d70701",
        1005 => x"3367b700",
        1006 => x"637ad700",
        1007 => x"3307e800",
        1008 => x"63660701",
        1009 => x"6374d700",
        1010 => x"33070701",
        1011 => x"3307d740",
        1012 => x"b356c702",
        1013 => x"3377c702",
        1014 => x"b386a602",
        1015 => x"93970701",
        1016 => x"13170701",
        1017 => x"93d70701",
        1018 => x"b3e7e700",
        1019 => x"63fad700",
        1020 => x"b307f800",
        1021 => x"63e60701",
        1022 => x"63f4d700",
        1023 => x"b3870701",
        1024 => x"b387d740",
        1025 => x"33d51701",
        1026 => x"93050000",
        1027 => x"67800000",
        1028 => x"37030001",
        1029 => x"93060001",
        1030 => x"e36666f4",
        1031 => x"93068001",
        1032 => x"6ff05ff4",
        1033 => x"93060000",
        1034 => x"630c0600",
        1035 => x"37070100",
        1036 => x"637ee606",
        1037 => x"93360610",
        1038 => x"93c61600",
        1039 => x"93963600",
        1040 => x"3357d600",
        1041 => x"b388e800",
        1042 => x"03c70800",
        1043 => x"3307d700",
        1044 => x"93060002",
        1045 => x"b388e640",
        1046 => x"6394e606",
        1047 => x"3387c540",
        1048 => x"93550801",
        1049 => x"3356b702",
        1050 => x"13150801",
        1051 => x"13550501",
        1052 => x"93d60701",
        1053 => x"3377b702",
        1054 => x"3306a602",
        1055 => x"13170701",
        1056 => x"33e7e600",
        1057 => x"637ac700",
        1058 => x"3307e800",
        1059 => x"63660701",
        1060 => x"6374c700",
        1061 => x"33070701",
        1062 => x"3307c740",
        1063 => x"b356b702",
        1064 => x"3377b702",
        1065 => x"b386a602",
        1066 => x"6ff05ff3",
        1067 => x"37070001",
        1068 => x"93060001",
        1069 => x"e366e6f8",
        1070 => x"93068001",
        1071 => x"6ff05ff8",
        1072 => x"33181601",
        1073 => x"b3d6e500",
        1074 => x"b3171501",
        1075 => x"b3951501",
        1076 => x"3357e500",
        1077 => x"13550801",
        1078 => x"3367b700",
        1079 => x"b3d5a602",
        1080 => x"13130801",
        1081 => x"13530301",
        1082 => x"b3f6a602",
        1083 => x"b3856502",
        1084 => x"13960601",
        1085 => x"93560701",
        1086 => x"b3e6c600",
        1087 => x"63fab600",
        1088 => x"b306d800",
        1089 => x"63e60601",
        1090 => x"63f4b600",
        1091 => x"b3860601",
        1092 => x"b386b640",
        1093 => x"33d6a602",
        1094 => x"13170701",
        1095 => x"13570701",
        1096 => x"b3f6a602",
        1097 => x"33066602",
        1098 => x"93960601",
        1099 => x"3367d700",
        1100 => x"637ac700",
        1101 => x"3307e800",
        1102 => x"63660701",
        1103 => x"6374c700",
        1104 => x"33070701",
        1105 => x"3307c740",
        1106 => x"6ff09ff1",
        1107 => x"63e4d51c",
        1108 => x"37080100",
        1109 => x"63fe0605",
        1110 => x"13b80610",
        1111 => x"13481800",
        1112 => x"13183800",
        1113 => x"b7380000",
        1114 => x"33d30601",
        1115 => x"938888d7",
        1116 => x"b3886800",
        1117 => x"83c80800",
        1118 => x"13030002",
        1119 => x"b3880801",
        1120 => x"33081341",
        1121 => x"63101305",
        1122 => x"63e4b600",
        1123 => x"636cc500",
        1124 => x"3306c540",
        1125 => x"b386d540",
        1126 => x"3337c500",
        1127 => x"93070600",
        1128 => x"3387e640",
        1129 => x"13850700",
        1130 => x"93050700",
        1131 => x"67800000",
        1132 => x"b7080001",
        1133 => x"13080001",
        1134 => x"e3e616fb",
        1135 => x"13088001",
        1136 => x"6ff05ffa",
        1137 => x"b3571601",
        1138 => x"b3960601",
        1139 => x"b3e6d700",
        1140 => x"33d71501",
        1141 => x"13de0601",
        1142 => x"335fc703",
        1143 => x"13930601",
        1144 => x"13530301",
        1145 => x"b3970501",
        1146 => x"b3551501",
        1147 => x"b3e5f500",
        1148 => x"93d70501",
        1149 => x"33160601",
        1150 => x"33150501",
        1151 => x"3377c703",
        1152 => x"b30ee303",
        1153 => x"13170701",
        1154 => x"b3e7e700",
        1155 => x"13070f00",
        1156 => x"63fed701",
        1157 => x"b387f600",
        1158 => x"1307ffff",
        1159 => x"63e8d700",
        1160 => x"63f6d701",
        1161 => x"1307efff",
        1162 => x"b387d700",
        1163 => x"b387d741",
        1164 => x"b3dec703",
        1165 => x"93950501",
        1166 => x"93d50501",
        1167 => x"b3f7c703",
        1168 => x"138e0e00",
        1169 => x"3303d303",
        1170 => x"93970701",
        1171 => x"b3e5f500",
        1172 => x"63fe6500",
        1173 => x"b385b600",
        1174 => x"138efeff",
        1175 => x"63e8d500",
        1176 => x"63f66500",
        1177 => x"138eeeff",
        1178 => x"b385d500",
        1179 => x"93170701",
        1180 => x"370f0100",
        1181 => x"b3e7c701",
        1182 => x"b3856540",
        1183 => x"1303ffff",
        1184 => x"33f76700",
        1185 => x"135e0601",
        1186 => x"93d70701",
        1187 => x"33736600",
        1188 => x"b30e6702",
        1189 => x"33836702",
        1190 => x"3307c703",
        1191 => x"b387c703",
        1192 => x"330e6700",
        1193 => x"13d70e01",
        1194 => x"3307c701",
        1195 => x"63746700",
        1196 => x"b387e701",
        1197 => x"13530701",
        1198 => x"b307f300",
        1199 => x"37030100",
        1200 => x"1303f3ff",
        1201 => x"33776700",
        1202 => x"13170701",
        1203 => x"b3fe6e00",
        1204 => x"3307d701",
        1205 => x"63e6f500",
        1206 => x"639ef500",
        1207 => x"637ce500",
        1208 => x"3306c740",
        1209 => x"3333c700",
        1210 => x"b306d300",
        1211 => x"13070600",
        1212 => x"b387d740",
        1213 => x"3307e540",
        1214 => x"3335e500",
        1215 => x"b385f540",
        1216 => x"b385a540",
        1217 => x"b3981501",
        1218 => x"33570701",
        1219 => x"33e5e800",
        1220 => x"b3d50501",
        1221 => x"67800000",
        1222 => x"13030500",
        1223 => x"630e0600",
        1224 => x"83830500",
        1225 => x"23007300",
        1226 => x"1306f6ff",
        1227 => x"13031300",
        1228 => x"93851500",
        1229 => x"e31606fe",
        1230 => x"67800000",
        1231 => x"13030500",
        1232 => x"630a0600",
        1233 => x"2300b300",
        1234 => x"1306f6ff",
        1235 => x"13031300",
        1236 => x"e31a06fe",
        1237 => x"67800000",
        1238 => x"630c0602",
        1239 => x"13030500",
        1240 => x"93061000",
        1241 => x"636ab500",
        1242 => x"9306f0ff",
        1243 => x"1307f6ff",
        1244 => x"3303e300",
        1245 => x"b385e500",
        1246 => x"83830500",
        1247 => x"23007300",
        1248 => x"1306f6ff",
        1249 => x"3303d300",
        1250 => x"b385d500",
        1251 => x"e31606fe",
        1252 => x"67800000",
        1253 => x"6f000000",
        1254 => x"130101ff",
        1255 => x"23248100",
        1256 => x"13040000",
        1257 => x"23229100",
        1258 => x"23202101",
        1259 => x"23261100",
        1260 => x"93040500",
        1261 => x"13090400",
        1262 => x"93070400",
        1263 => x"732410c8",
        1264 => x"732910c0",
        1265 => x"f32710c8",
        1266 => x"e31af4fe",
        1267 => x"37460f00",
        1268 => x"13060624",
        1269 => x"93060000",
        1270 => x"13050900",
        1271 => x"93050400",
        1272 => x"eff05fb5",
        1273 => x"37460f00",
        1274 => x"23a4a400",
        1275 => x"93050400",
        1276 => x"13050900",
        1277 => x"13060624",
        1278 => x"93060000",
        1279 => x"eff08ff0",
        1280 => x"8320c100",
        1281 => x"03248100",
        1282 => x"23a0a400",
        1283 => x"23a2b400",
        1284 => x"03290100",
        1285 => x"83244100",
        1286 => x"13050000",
        1287 => x"13010101",
        1288 => x"67800000",
        1289 => x"03a74188",
        1290 => x"b7870020",
        1291 => x"93870700",
        1292 => x"93060040",
        1293 => x"b387d740",
        1294 => x"630c0700",
        1295 => x"3305a700",
        1296 => x"63e2a702",
        1297 => x"23a2a188",
        1298 => x"13050700",
        1299 => x"67800000",
        1300 => x"93868189",
        1301 => x"13878189",
        1302 => x"23a2d188",
        1303 => x"3305a700",
        1304 => x"e3f2a7fe",
        1305 => x"130101ff",
        1306 => x"23261100",
        1307 => x"ef00403d",
        1308 => x"8320c100",
        1309 => x"9307c000",
        1310 => x"2320f500",
        1311 => x"1307f0ff",
        1312 => x"13050700",
        1313 => x"13010101",
        1314 => x"67800000",
        1315 => x"370700f0",
        1316 => x"83274702",
        1317 => x"93f74700",
        1318 => x"e38c07fe",
        1319 => x"03258702",
        1320 => x"1375f50f",
        1321 => x"67800000",
        1322 => x"f32710fc",
        1323 => x"63960700",
        1324 => x"b7f7fa02",
        1325 => x"93870708",
        1326 => x"63060500",
        1327 => x"33d5a702",
        1328 => x"1305f5ff",
        1329 => x"b70700f0",
        1330 => x"23a6a702",
        1331 => x"23a0b702",
        1332 => x"67800000",
        1333 => x"1375f50f",
        1334 => x"b70700f0",
        1335 => x"370700f0",
        1336 => x"23a4a702",
        1337 => x"83274702",
        1338 => x"93f70701",
        1339 => x"e38c07fe",
        1340 => x"67800000",
        1341 => x"630e0502",
        1342 => x"130101ff",
        1343 => x"23248100",
        1344 => x"23261100",
        1345 => x"13040500",
        1346 => x"03450500",
        1347 => x"630a0500",
        1348 => x"13041400",
        1349 => x"eff01ffc",
        1350 => x"03450400",
        1351 => x"e31a05fe",
        1352 => x"8320c100",
        1353 => x"03248100",
        1354 => x"13010101",
        1355 => x"67800000",
        1356 => x"67800000",
        1357 => x"130101f9",
        1358 => x"23248106",
        1359 => x"23229106",
        1360 => x"23261106",
        1361 => x"23202107",
        1362 => x"232e3105",
        1363 => x"232c4105",
        1364 => x"232a5105",
        1365 => x"23286105",
        1366 => x"23267105",
        1367 => x"23248105",
        1368 => x"23229105",
        1369 => x"2320a105",
        1370 => x"93040500",
        1371 => x"13840500",
        1372 => x"232c0100",
        1373 => x"232e0100",
        1374 => x"23200102",
        1375 => x"23220102",
        1376 => x"23240102",
        1377 => x"23260102",
        1378 => x"23280102",
        1379 => x"232a0102",
        1380 => x"232c0102",
        1381 => x"232e0102",
        1382 => x"97f2ffff",
        1383 => x"9382c2cf",
        1384 => x"73905230",
        1385 => x"37c50100",
        1386 => x"93050004",
        1387 => x"13050520",
        1388 => x"eff09fef",
        1389 => x"37877d01",
        1390 => x"b70700f0",
        1391 => x"1307f783",
        1392 => x"23a6e708",
        1393 => x"93061001",
        1394 => x"37170000",
        1395 => x"23a0d708",
        1396 => x"13077738",
        1397 => x"23a8e70a",
        1398 => x"37270000",
        1399 => x"1307f770",
        1400 => x"23a6e70a",
        1401 => x"23a0d70a",
        1402 => x"13078070",
        1403 => x"23a0e706",
        1404 => x"3707f900",
        1405 => x"13078700",
        1406 => x"23a0e704",
        1407 => x"1307a007",
        1408 => x"23ace700",
        1409 => x"93020008",
        1410 => x"73904230",
        1411 => x"b7220000",
        1412 => x"93828280",
        1413 => x"73900230",
        1414 => x"b7390000",
        1415 => x"138549ec",
        1416 => x"eff05fed",
        1417 => x"63549002",
        1418 => x"1389f4ff",
        1419 => x"9304f0ff",
        1420 => x"03250400",
        1421 => x"1309f9ff",
        1422 => x"13044400",
        1423 => x"eff09feb",
        1424 => x"138549ec",
        1425 => x"eff01feb",
        1426 => x"e31499fe",
        1427 => x"37350000",
        1428 => x"b7faeeee",
        1429 => x"130585e9",
        1430 => x"b7090010",
        1431 => x"37140000",
        1432 => x"1389faee",
        1433 => x"eff01fe9",
        1434 => x"373b0000",
        1435 => x"9389f9ff",
        1436 => x"938aeaee",
        1437 => x"130404e1",
        1438 => x"93040000",
        1439 => x"b71b0000",
        1440 => x"938b0b2c",
        1441 => x"130af000",
        1442 => x"93050000",
        1443 => x"13058100",
        1444 => x"ef008036",
        1445 => x"938bfbff",
        1446 => x"630a0502",
        1447 => x"e3960bfe",
        1448 => x"73001000",
        1449 => x"b70700f0",
        1450 => x"9306f00f",
        1451 => x"23a4d706",
        1452 => x"03a70704",
        1453 => x"93860704",
        1454 => x"13670730",
        1455 => x"23a0e704",
        1456 => x"93070009",
        1457 => x"23a4f600",
        1458 => x"6ff05ffb",
        1459 => x"032c8100",
        1460 => x"8325c100",
        1461 => x"13060400",
        1462 => x"9357cc01",
        1463 => x"13974500",
        1464 => x"b367f700",
        1465 => x"b3f73701",
        1466 => x"33773c01",
        1467 => x"13d5f541",
        1468 => x"13d88501",
        1469 => x"3307f700",
        1470 => x"33070701",
        1471 => x"9377d500",
        1472 => x"3307f700",
        1473 => x"33774703",
        1474 => x"937725ff",
        1475 => x"93860400",
        1476 => x"13050c00",
        1477 => x"3307f700",
        1478 => x"b307ec40",
        1479 => x"1357f741",
        1480 => x"3338fc00",
        1481 => x"3387e540",
        1482 => x"33070741",
        1483 => x"b3885703",
        1484 => x"33072703",
        1485 => x"33b82703",
        1486 => x"33071701",
        1487 => x"b3872703",
        1488 => x"33070701",
        1489 => x"1358f741",
        1490 => x"13783800",
        1491 => x"b307f800",
        1492 => x"33b80701",
        1493 => x"3307e800",
        1494 => x"1318e701",
        1495 => x"93d72700",
        1496 => x"b367f800",
        1497 => x"13582740",
        1498 => x"93184800",
        1499 => x"13d3c701",
        1500 => x"33e36800",
        1501 => x"33733301",
        1502 => x"b3f83701",
        1503 => x"135e8801",
        1504 => x"1357f741",
        1505 => x"b3886800",
        1506 => x"b388c801",
        1507 => x"1373d700",
        1508 => x"b3886800",
        1509 => x"b3f84803",
        1510 => x"137727ff",
        1511 => x"939c4700",
        1512 => x"b38cfc40",
        1513 => x"939c2c00",
        1514 => x"b30c9c41",
        1515 => x"b388e800",
        1516 => x"33871741",
        1517 => x"93d8f841",
        1518 => x"33b3e700",
        1519 => x"33081841",
        1520 => x"33086840",
        1521 => x"33082803",
        1522 => x"33035703",
        1523 => x"b3382703",
        1524 => x"33086800",
        1525 => x"33072703",
        1526 => x"33081801",
        1527 => x"9358f841",
        1528 => x"93f83800",
        1529 => x"3387e800",
        1530 => x"b3381701",
        1531 => x"b3880801",
        1532 => x"9398e801",
        1533 => x"13572700",
        1534 => x"33e7e800",
        1535 => x"13184700",
        1536 => x"3307e840",
        1537 => x"13172700",
        1538 => x"338de740",
        1539 => x"efe01fe8",
        1540 => x"83260101",
        1541 => x"13070500",
        1542 => x"13880c00",
        1543 => x"93070d00",
        1544 => x"13060c00",
        1545 => x"93058bec",
        1546 => x"13058101",
        1547 => x"ef00c015",
        1548 => x"13058101",
        1549 => x"eff01fcc",
        1550 => x"e3980be4",
        1551 => x"6ff05fe6",
        1552 => x"03a5c187",
        1553 => x"67800000",
        1554 => x"130101ff",
        1555 => x"23248100",
        1556 => x"23261100",
        1557 => x"93070000",
        1558 => x"13040500",
        1559 => x"63880700",
        1560 => x"93050000",
        1561 => x"97000000",
        1562 => x"e7000000",
        1563 => x"b7370000",
        1564 => x"03a58702",
        1565 => x"83278502",
        1566 => x"63840700",
        1567 => x"e7800700",
        1568 => x"13050400",
        1569 => x"eff01fb1",
        1570 => x"130101ff",
        1571 => x"23248100",
        1572 => x"23229100",
        1573 => x"37340000",
        1574 => x"b7340000",
        1575 => x"9387c402",
        1576 => x"1304c402",
        1577 => x"3304f440",
        1578 => x"23202101",
        1579 => x"23261100",
        1580 => x"13542440",
        1581 => x"9384c402",
        1582 => x"13090000",
        1583 => x"63108904",
        1584 => x"b7340000",
        1585 => x"37340000",
        1586 => x"9387c402",
        1587 => x"1304c402",
        1588 => x"3304f440",
        1589 => x"13542440",
        1590 => x"9384c402",
        1591 => x"13090000",
        1592 => x"63188902",
        1593 => x"8320c100",
        1594 => x"03248100",
        1595 => x"83244100",
        1596 => x"03290100",
        1597 => x"13010101",
        1598 => x"67800000",
        1599 => x"83a70400",
        1600 => x"13091900",
        1601 => x"93844400",
        1602 => x"e7800700",
        1603 => x"6ff01ffb",
        1604 => x"83a70400",
        1605 => x"13091900",
        1606 => x"93844400",
        1607 => x"e7800700",
        1608 => x"6ff01ffc",
        1609 => x"130101f6",
        1610 => x"232af108",
        1611 => x"b7070080",
        1612 => x"93c7f7ff",
        1613 => x"232ef100",
        1614 => x"2328f100",
        1615 => x"b707ffff",
        1616 => x"2326d108",
        1617 => x"2324b100",
        1618 => x"232cb100",
        1619 => x"93878720",
        1620 => x"9306c108",
        1621 => x"93058100",
        1622 => x"232e1106",
        1623 => x"232af100",
        1624 => x"2328e108",
        1625 => x"232c0109",
        1626 => x"232e1109",
        1627 => x"2322d100",
        1628 => x"ef00c040",
        1629 => x"83278100",
        1630 => x"23800700",
        1631 => x"8320c107",
        1632 => x"1301010a",
        1633 => x"67800000",
        1634 => x"130101f6",
        1635 => x"232af108",
        1636 => x"b7070080",
        1637 => x"93c7f7ff",
        1638 => x"232ef100",
        1639 => x"2328f100",
        1640 => x"b707ffff",
        1641 => x"93878720",
        1642 => x"232af100",
        1643 => x"2324a100",
        1644 => x"232ca100",
        1645 => x"03a5c187",
        1646 => x"2324c108",
        1647 => x"2326d108",
        1648 => x"13860500",
        1649 => x"93068108",
        1650 => x"93058100",
        1651 => x"232e1106",
        1652 => x"2328e108",
        1653 => x"232c0109",
        1654 => x"232e1109",
        1655 => x"2322d100",
        1656 => x"ef00c039",
        1657 => x"83278100",
        1658 => x"23800700",
        1659 => x"8320c107",
        1660 => x"1301010a",
        1661 => x"67800000",
        1662 => x"13860500",
        1663 => x"93050500",
        1664 => x"03a5c187",
        1665 => x"6f004000",
        1666 => x"130101ff",
        1667 => x"23248100",
        1668 => x"23229100",
        1669 => x"13040500",
        1670 => x"13850500",
        1671 => x"93050600",
        1672 => x"23261100",
        1673 => x"23a40188",
        1674 => x"eff01f97",
        1675 => x"9307f0ff",
        1676 => x"6318f500",
        1677 => x"83a78188",
        1678 => x"63840700",
        1679 => x"2320f400",
        1680 => x"8320c100",
        1681 => x"03248100",
        1682 => x"83244100",
        1683 => x"13010101",
        1684 => x"67800000",
        1685 => x"130101fe",
        1686 => x"23282101",
        1687 => x"03a98500",
        1688 => x"232c8100",
        1689 => x"23263101",
        1690 => x"23225101",
        1691 => x"23206101",
        1692 => x"232e1100",
        1693 => x"232a9100",
        1694 => x"23244101",
        1695 => x"83aa0500",
        1696 => x"13840500",
        1697 => x"130b0600",
        1698 => x"93890600",
        1699 => x"63ec2609",
        1700 => x"8397c500",
        1701 => x"13f70748",
        1702 => x"63040708",
        1703 => x"03274401",
        1704 => x"93043000",
        1705 => x"83a50501",
        1706 => x"b384e402",
        1707 => x"13072000",
        1708 => x"b38aba40",
        1709 => x"130a0500",
        1710 => x"b3c4e402",
        1711 => x"13871600",
        1712 => x"33075701",
        1713 => x"63f4e400",
        1714 => x"93040700",
        1715 => x"93f70740",
        1716 => x"6386070a",
        1717 => x"93850400",
        1718 => x"13050a00",
        1719 => x"ef001067",
        1720 => x"13090500",
        1721 => x"630c050a",
        1722 => x"83250401",
        1723 => x"13860a00",
        1724 => x"eff09f82",
        1725 => x"8357c400",
        1726 => x"93f7f7b7",
        1727 => x"93e70708",
        1728 => x"2316f400",
        1729 => x"23282401",
        1730 => x"232a9400",
        1731 => x"33095901",
        1732 => x"b3845441",
        1733 => x"23202401",
        1734 => x"23249400",
        1735 => x"13890900",
        1736 => x"63f42901",
        1737 => x"13890900",
        1738 => x"03250400",
        1739 => x"13060900",
        1740 => x"93050b00",
        1741 => x"eff05f82",
        1742 => x"83278400",
        1743 => x"13050000",
        1744 => x"b3872741",
        1745 => x"2324f400",
        1746 => x"83270400",
        1747 => x"b3872701",
        1748 => x"2320f400",
        1749 => x"8320c101",
        1750 => x"03248101",
        1751 => x"83244101",
        1752 => x"03290101",
        1753 => x"8329c100",
        1754 => x"032a8100",
        1755 => x"832a4100",
        1756 => x"032b0100",
        1757 => x"13010102",
        1758 => x"67800000",
        1759 => x"13860400",
        1760 => x"13050a00",
        1761 => x"ef001071",
        1762 => x"13090500",
        1763 => x"e31c05f6",
        1764 => x"83250401",
        1765 => x"13050a00",
        1766 => x"ef00d04b",
        1767 => x"9307c000",
        1768 => x"2320fa00",
        1769 => x"8357c400",
        1770 => x"1305f0ff",
        1771 => x"93e70704",
        1772 => x"2316f400",
        1773 => x"6ff01ffa",
        1774 => x"83278600",
        1775 => x"130101fd",
        1776 => x"232e3101",
        1777 => x"23286101",
        1778 => x"23261102",
        1779 => x"23248102",
        1780 => x"23229102",
        1781 => x"23202103",
        1782 => x"232c4101",
        1783 => x"232a5101",
        1784 => x"23267101",
        1785 => x"23248101",
        1786 => x"23229101",
        1787 => x"2320a101",
        1788 => x"032b0600",
        1789 => x"93090600",
        1790 => x"63940712",
        1791 => x"13050000",
        1792 => x"8320c102",
        1793 => x"03248102",
        1794 => x"23a20900",
        1795 => x"83244102",
        1796 => x"03290102",
        1797 => x"8329c101",
        1798 => x"032a8101",
        1799 => x"832a4101",
        1800 => x"032b0101",
        1801 => x"832bc100",
        1802 => x"032c8100",
        1803 => x"832c4100",
        1804 => x"032d0100",
        1805 => x"13010103",
        1806 => x"67800000",
        1807 => x"832b0b00",
        1808 => x"032d4b00",
        1809 => x"130b8b00",
        1810 => x"03298400",
        1811 => x"832a0400",
        1812 => x"e3060dfe",
        1813 => x"63642d09",
        1814 => x"8317c400",
        1815 => x"13f70748",
        1816 => x"630e0706",
        1817 => x"83244401",
        1818 => x"83250401",
        1819 => x"b3049c02",
        1820 => x"b38aba40",
        1821 => x"13871a00",
        1822 => x"3307a701",
        1823 => x"b3c49403",
        1824 => x"63f4e400",
        1825 => x"93040700",
        1826 => x"93f70740",
        1827 => x"6388070a",
        1828 => x"93850400",
        1829 => x"13050a00",
        1830 => x"ef00504b",
        1831 => x"13090500",
        1832 => x"630e050a",
        1833 => x"83250401",
        1834 => x"13860a00",
        1835 => x"eff0cfe6",
        1836 => x"8357c400",
        1837 => x"93f7f7b7",
        1838 => x"93e70708",
        1839 => x"2316f400",
        1840 => x"23282401",
        1841 => x"232a9400",
        1842 => x"33095901",
        1843 => x"b3845441",
        1844 => x"23202401",
        1845 => x"23249400",
        1846 => x"13090d00",
        1847 => x"63742d01",
        1848 => x"13090d00",
        1849 => x"03250400",
        1850 => x"13060900",
        1851 => x"93850b00",
        1852 => x"eff08fe6",
        1853 => x"83278400",
        1854 => x"b3872741",
        1855 => x"2324f400",
        1856 => x"83270400",
        1857 => x"b3872701",
        1858 => x"2320f400",
        1859 => x"83a78900",
        1860 => x"b387a741",
        1861 => x"23a4f900",
        1862 => x"e39207f2",
        1863 => x"6ff01fee",
        1864 => x"130a0500",
        1865 => x"13840500",
        1866 => x"930b0000",
        1867 => x"130d0000",
        1868 => x"130c3000",
        1869 => x"930c2000",
        1870 => x"6ff01ff1",
        1871 => x"13860400",
        1872 => x"13050a00",
        1873 => x"ef001055",
        1874 => x"13090500",
        1875 => x"e31a05f6",
        1876 => x"83250401",
        1877 => x"13050a00",
        1878 => x"ef00d02f",
        1879 => x"9307c000",
        1880 => x"2320fa00",
        1881 => x"8357c400",
        1882 => x"1305f0ff",
        1883 => x"93e70704",
        1884 => x"2316f400",
        1885 => x"23a40900",
        1886 => x"6ff09fe8",
        1887 => x"83d7c500",
        1888 => x"130101f5",
        1889 => x"2324810a",
        1890 => x"2322910a",
        1891 => x"2320210b",
        1892 => x"232c4109",
        1893 => x"2326110a",
        1894 => x"232e3109",
        1895 => x"232a5109",
        1896 => x"23286109",
        1897 => x"23267109",
        1898 => x"23248109",
        1899 => x"23229109",
        1900 => x"2320a109",
        1901 => x"232eb107",
        1902 => x"93f70708",
        1903 => x"130a0500",
        1904 => x"13890500",
        1905 => x"93040600",
        1906 => x"13840600",
        1907 => x"63880706",
        1908 => x"83a70501",
        1909 => x"63940706",
        1910 => x"93050004",
        1911 => x"ef001037",
        1912 => x"2320a900",
        1913 => x"2328a900",
        1914 => x"63160504",
        1915 => x"9307c000",
        1916 => x"2320fa00",
        1917 => x"1305f0ff",
        1918 => x"8320c10a",
        1919 => x"0324810a",
        1920 => x"8324410a",
        1921 => x"0329010a",
        1922 => x"8329c109",
        1923 => x"032a8109",
        1924 => x"832a4109",
        1925 => x"032b0109",
        1926 => x"832bc108",
        1927 => x"032c8108",
        1928 => x"832c4108",
        1929 => x"032d0108",
        1930 => x"832dc107",
        1931 => x"1301010b",
        1932 => x"67800000",
        1933 => x"93070004",
        1934 => x"232af900",
        1935 => x"93070002",
        1936 => x"a304f102",
        1937 => x"93070003",
        1938 => x"23220102",
        1939 => x"2305f102",
        1940 => x"23268100",
        1941 => x"930c5002",
        1942 => x"373b0000",
        1943 => x"b73b0000",
        1944 => x"373d0000",
        1945 => x"372c0000",
        1946 => x"930a0000",
        1947 => x"13840400",
        1948 => x"83470400",
        1949 => x"63840700",
        1950 => x"639c970d",
        1951 => x"b30d9440",
        1952 => x"63069402",
        1953 => x"93860d00",
        1954 => x"13860400",
        1955 => x"93050900",
        1956 => x"13050a00",
        1957 => x"eff01fbc",
        1958 => x"9307f0ff",
        1959 => x"6304f524",
        1960 => x"83274102",
        1961 => x"b387b701",
        1962 => x"2322f102",
        1963 => x"83470400",
        1964 => x"638a0722",
        1965 => x"9307f0ff",
        1966 => x"93041400",
        1967 => x"23280100",
        1968 => x"232e0100",
        1969 => x"232af100",
        1970 => x"232c0100",
        1971 => x"a3090104",
        1972 => x"23240106",
        1973 => x"930d1000",
        1974 => x"83c50400",
        1975 => x"13065000",
        1976 => x"13054bf9",
        1977 => x"ef00d014",
        1978 => x"83270101",
        1979 => x"13841400",
        1980 => x"63140506",
        1981 => x"13f70701",
        1982 => x"63060700",
        1983 => x"13070002",
        1984 => x"a309e104",
        1985 => x"13f78700",
        1986 => x"63060700",
        1987 => x"1307b002",
        1988 => x"a309e104",
        1989 => x"83c60400",
        1990 => x"1307a002",
        1991 => x"638ce604",
        1992 => x"8327c101",
        1993 => x"13840400",
        1994 => x"93060000",
        1995 => x"13069000",
        1996 => x"1305a000",
        1997 => x"03470400",
        1998 => x"93051400",
        1999 => x"130707fd",
        2000 => x"637ee608",
        2001 => x"63840604",
        2002 => x"232ef100",
        2003 => x"6f000004",
        2004 => x"13041400",
        2005 => x"6ff0dff1",
        2006 => x"13074bf9",
        2007 => x"3305e540",
        2008 => x"3395ad00",
        2009 => x"b3e7a700",
        2010 => x"2328f100",
        2011 => x"93040400",
        2012 => x"6ff09ff6",
        2013 => x"0327c100",
        2014 => x"93064700",
        2015 => x"03270700",
        2016 => x"2326d100",
        2017 => x"63420704",
        2018 => x"232ee100",
        2019 => x"03470400",
        2020 => x"9307e002",
        2021 => x"6314f708",
        2022 => x"03471400",
        2023 => x"9307a002",
        2024 => x"6318f704",
        2025 => x"8327c100",
        2026 => x"13042400",
        2027 => x"13874700",
        2028 => x"83a70700",
        2029 => x"2326e100",
        2030 => x"63d40700",
        2031 => x"9307f0ff",
        2032 => x"232af100",
        2033 => x"6f008005",
        2034 => x"3307e040",
        2035 => x"93e72700",
        2036 => x"232ee100",
        2037 => x"2328f100",
        2038 => x"6ff05ffb",
        2039 => x"b387a702",
        2040 => x"13840500",
        2041 => x"93061000",
        2042 => x"b387e700",
        2043 => x"6ff09ff4",
        2044 => x"13041400",
        2045 => x"232a0100",
        2046 => x"93060000",
        2047 => x"93070000",
        2048 => x"13069000",
        2049 => x"1305a000",
        2050 => x"03470400",
        2051 => x"93051400",
        2052 => x"130707fd",
        2053 => x"6372e608",
        2054 => x"e39406fa",
        2055 => x"83450400",
        2056 => x"13063000",
        2057 => x"1385cbf9",
        2058 => x"ef009000",
        2059 => x"63020502",
        2060 => x"9387cbf9",
        2061 => x"3305f540",
        2062 => x"83270101",
        2063 => x"13070004",
        2064 => x"3317a700",
        2065 => x"b3e7e700",
        2066 => x"13041400",
        2067 => x"2328f100",
        2068 => x"83450400",
        2069 => x"13066000",
        2070 => x"13050dfa",
        2071 => x"93041400",
        2072 => x"2304b102",
        2073 => x"ef00c07c",
        2074 => x"63080508",
        2075 => x"63980a04",
        2076 => x"03270101",
        2077 => x"8327c100",
        2078 => x"13770710",
        2079 => x"63080702",
        2080 => x"93874700",
        2081 => x"2326f100",
        2082 => x"83274102",
        2083 => x"b3873701",
        2084 => x"2322f102",
        2085 => x"6ff09fdd",
        2086 => x"b387a702",
        2087 => x"13840500",
        2088 => x"93061000",
        2089 => x"b387e700",
        2090 => x"6ff01ff6",
        2091 => x"93877700",
        2092 => x"93f787ff",
        2093 => x"93878700",
        2094 => x"6ff0dffc",
        2095 => x"1307c100",
        2096 => x"93064ca5",
        2097 => x"13060900",
        2098 => x"93050101",
        2099 => x"13050a00",
        2100 => x"97000000",
        2101 => x"e7000000",
        2102 => x"9307f0ff",
        2103 => x"93090500",
        2104 => x"e314f5fa",
        2105 => x"8357c900",
        2106 => x"93f70704",
        2107 => x"e39407d0",
        2108 => x"03254102",
        2109 => x"6ff05fd0",
        2110 => x"1307c100",
        2111 => x"93064ca5",
        2112 => x"13060900",
        2113 => x"93050101",
        2114 => x"13050a00",
        2115 => x"ef00801b",
        2116 => x"6ff09ffc",
        2117 => x"130101fd",
        2118 => x"232a5101",
        2119 => x"83a70501",
        2120 => x"930a0700",
        2121 => x"03a78500",
        2122 => x"23248102",
        2123 => x"23202103",
        2124 => x"232e3101",
        2125 => x"232c4101",
        2126 => x"23261102",
        2127 => x"23229102",
        2128 => x"23286101",
        2129 => x"23267101",
        2130 => x"93090500",
        2131 => x"13840500",
        2132 => x"13090600",
        2133 => x"138a0600",
        2134 => x"63d4e700",
        2135 => x"93070700",
        2136 => x"2320f900",
        2137 => x"03473404",
        2138 => x"63060700",
        2139 => x"93871700",
        2140 => x"2320f900",
        2141 => x"83270400",
        2142 => x"93f70702",
        2143 => x"63880700",
        2144 => x"83270900",
        2145 => x"93872700",
        2146 => x"2320f900",
        2147 => x"83240400",
        2148 => x"93f46400",
        2149 => x"639e0400",
        2150 => x"130b9401",
        2151 => x"930bf0ff",
        2152 => x"8327c400",
        2153 => x"03270900",
        2154 => x"b387e740",
        2155 => x"63c2f408",
        2156 => x"83473404",
        2157 => x"b336f000",
        2158 => x"83270400",
        2159 => x"93f70702",
        2160 => x"6390070c",
        2161 => x"13063404",
        2162 => x"93050a00",
        2163 => x"13850900",
        2164 => x"e7800a00",
        2165 => x"9307f0ff",
        2166 => x"6308f506",
        2167 => x"83270400",
        2168 => x"13074000",
        2169 => x"93040000",
        2170 => x"93f76700",
        2171 => x"639ce700",
        2172 => x"8324c400",
        2173 => x"83270900",
        2174 => x"b384f440",
        2175 => x"63d40400",
        2176 => x"93040000",
        2177 => x"83278400",
        2178 => x"03270401",
        2179 => x"6356f700",
        2180 => x"b387e740",
        2181 => x"b384f400",
        2182 => x"13090000",
        2183 => x"1304a401",
        2184 => x"130bf0ff",
        2185 => x"63902409",
        2186 => x"13050000",
        2187 => x"6f000002",
        2188 => x"93061000",
        2189 => x"13060b00",
        2190 => x"93050a00",
        2191 => x"13850900",
        2192 => x"e7800a00",
        2193 => x"631a7503",
        2194 => x"1305f0ff",
        2195 => x"8320c102",
        2196 => x"03248102",
        2197 => x"83244102",
        2198 => x"03290102",
        2199 => x"8329c101",
        2200 => x"032a8101",
        2201 => x"832a4101",
        2202 => x"032b0101",
        2203 => x"832bc100",
        2204 => x"13010103",
        2205 => x"67800000",
        2206 => x"93841400",
        2207 => x"6ff05ff2",
        2208 => x"3307d400",
        2209 => x"13060003",
        2210 => x"a301c704",
        2211 => x"03475404",
        2212 => x"93871600",
        2213 => x"b307f400",
        2214 => x"93862600",
        2215 => x"a381e704",
        2216 => x"6ff05ff2",
        2217 => x"93061000",
        2218 => x"13060400",
        2219 => x"93050a00",
        2220 => x"13850900",
        2221 => x"e7800a00",
        2222 => x"e30865f9",
        2223 => x"13091900",
        2224 => x"6ff05ff6",
        2225 => x"130101fd",
        2226 => x"23248102",
        2227 => x"23229102",
        2228 => x"23202103",
        2229 => x"232e3101",
        2230 => x"23261102",
        2231 => x"232c4101",
        2232 => x"232a5101",
        2233 => x"23286101",
        2234 => x"83c88501",
        2235 => x"93078007",
        2236 => x"93040500",
        2237 => x"13840500",
        2238 => x"13090600",
        2239 => x"93890600",
        2240 => x"63ee1701",
        2241 => x"93072006",
        2242 => x"93863504",
        2243 => x"63ee1701",
        2244 => x"638a082a",
        2245 => x"93078005",
        2246 => x"638af820",
        2247 => x"930a2404",
        2248 => x"23011405",
        2249 => x"6f004004",
        2250 => x"9387d8f9",
        2251 => x"93f7f70f",
        2252 => x"13065001",
        2253 => x"e364f6fe",
        2254 => x"37360000",
        2255 => x"93972700",
        2256 => x"130606fd",
        2257 => x"b387c700",
        2258 => x"83a70700",
        2259 => x"67800700",
        2260 => x"83270700",
        2261 => x"938a2504",
        2262 => x"93864700",
        2263 => x"83a70700",
        2264 => x"2320d700",
        2265 => x"2381f504",
        2266 => x"93071000",
        2267 => x"6f004029",
        2268 => x"03a60500",
        2269 => x"83270700",
        2270 => x"13750608",
        2271 => x"93854700",
        2272 => x"630e0504",
        2273 => x"83a70700",
        2274 => x"2320b700",
        2275 => x"37370000",
        2276 => x"83254400",
        2277 => x"130887fa",
        2278 => x"63d2071e",
        2279 => x"1307d002",
        2280 => x"a301e404",
        2281 => x"2324b400",
        2282 => x"63d80504",
        2283 => x"b307f040",
        2284 => x"1307a000",
        2285 => x"938a0600",
        2286 => x"33f6e702",
        2287 => x"938afaff",
        2288 => x"3306c800",
        2289 => x"03460600",
        2290 => x"2380ca00",
        2291 => x"13860700",
        2292 => x"b3d7e702",
        2293 => x"e372e6fe",
        2294 => x"6f008009",
        2295 => x"83a70700",
        2296 => x"13750604",
        2297 => x"2320b700",
        2298 => x"e30205fa",
        2299 => x"93970701",
        2300 => x"93d70741",
        2301 => x"6ff09ff9",
        2302 => x"1376b6ff",
        2303 => x"2320c400",
        2304 => x"6ff0dffa",
        2305 => x"03a60500",
        2306 => x"83270700",
        2307 => x"13750608",
        2308 => x"93854700",
        2309 => x"63080500",
        2310 => x"2320b700",
        2311 => x"83a70700",
        2312 => x"6f004001",
        2313 => x"13760604",
        2314 => x"2320b700",
        2315 => x"e30806fe",
        2316 => x"83d70700",
        2317 => x"37380000",
        2318 => x"1307f006",
        2319 => x"130888fa",
        2320 => x"639ae812",
        2321 => x"13078000",
        2322 => x"a3010404",
        2323 => x"03264400",
        2324 => x"2324c400",
        2325 => x"e34006f6",
        2326 => x"83250400",
        2327 => x"93f5b5ff",
        2328 => x"2320b400",
        2329 => x"e39807f4",
        2330 => x"938a0600",
        2331 => x"e31406f4",
        2332 => x"93078000",
        2333 => x"6314f702",
        2334 => x"83270400",
        2335 => x"93f71700",
        2336 => x"638e0700",
        2337 => x"03274400",
        2338 => x"83270401",
        2339 => x"63c8e700",
        2340 => x"93070003",
        2341 => x"a38ffafe",
        2342 => x"938afaff",
        2343 => x"b3865641",
        2344 => x"2328d400",
        2345 => x"13870900",
        2346 => x"93060900",
        2347 => x"1306c100",
        2348 => x"93050400",
        2349 => x"13850400",
        2350 => x"eff0dfc5",
        2351 => x"130af0ff",
        2352 => x"63164515",
        2353 => x"1305f0ff",
        2354 => x"8320c102",
        2355 => x"03248102",
        2356 => x"83244102",
        2357 => x"03290102",
        2358 => x"8329c101",
        2359 => x"032a8101",
        2360 => x"832a4101",
        2361 => x"032b0101",
        2362 => x"13010103",
        2363 => x"67800000",
        2364 => x"83a70500",
        2365 => x"93e70702",
        2366 => x"23a0f500",
        2367 => x"37380000",
        2368 => x"93088007",
        2369 => x"1308c8fb",
        2370 => x"03260400",
        2371 => x"a3021405",
        2372 => x"83270700",
        2373 => x"13750608",
        2374 => x"93854700",
        2375 => x"630e0500",
        2376 => x"2320b700",
        2377 => x"83a70700",
        2378 => x"6f000002",
        2379 => x"37380000",
        2380 => x"130888fa",
        2381 => x"6ff05ffd",
        2382 => x"13750604",
        2383 => x"2320b700",
        2384 => x"e30205fe",
        2385 => x"83d70700",
        2386 => x"13771600",
        2387 => x"63060700",
        2388 => x"13660602",
        2389 => x"2320c400",
        2390 => x"63860700",
        2391 => x"13070001",
        2392 => x"6ff09fee",
        2393 => x"03270400",
        2394 => x"1377f7fd",
        2395 => x"2320e400",
        2396 => x"6ff0dffe",
        2397 => x"1307a000",
        2398 => x"6ff01fed",
        2399 => x"130887fa",
        2400 => x"1307a000",
        2401 => x"6ff09fec",
        2402 => x"03a60500",
        2403 => x"83270700",
        2404 => x"83a54501",
        2405 => x"13780608",
        2406 => x"13854700",
        2407 => x"630a0800",
        2408 => x"2320a700",
        2409 => x"83a70700",
        2410 => x"23a0b700",
        2411 => x"6f008001",
        2412 => x"2320a700",
        2413 => x"13760604",
        2414 => x"83a70700",
        2415 => x"e30606fe",
        2416 => x"2390b700",
        2417 => x"23280400",
        2418 => x"938a0600",
        2419 => x"6ff09fed",
        2420 => x"83270700",
        2421 => x"03a64500",
        2422 => x"93050000",
        2423 => x"93864700",
        2424 => x"2320d700",
        2425 => x"83aa0700",
        2426 => x"13850a00",
        2427 => x"ef004024",
        2428 => x"63060500",
        2429 => x"33055541",
        2430 => x"2322a400",
        2431 => x"83274400",
        2432 => x"2328f400",
        2433 => x"a3010404",
        2434 => x"6ff0dfe9",
        2435 => x"83260401",
        2436 => x"13860a00",
        2437 => x"93050900",
        2438 => x"13850400",
        2439 => x"e7800900",
        2440 => x"e30245eb",
        2441 => x"83270400",
        2442 => x"93f72700",
        2443 => x"63940704",
        2444 => x"8327c100",
        2445 => x"0325c400",
        2446 => x"e358f5e8",
        2447 => x"13850700",
        2448 => x"6ff09fe8",
        2449 => x"93061000",
        2450 => x"13860a00",
        2451 => x"93050900",
        2452 => x"13850400",
        2453 => x"e7800900",
        2454 => x"e30665e7",
        2455 => x"130a1a00",
        2456 => x"8327c400",
        2457 => x"0327c100",
        2458 => x"b387e740",
        2459 => x"e34cfafc",
        2460 => x"6ff01ffc",
        2461 => x"130a0000",
        2462 => x"930a9401",
        2463 => x"130bf0ff",
        2464 => x"6ff01ffe",
        2465 => x"130101ff",
        2466 => x"23248100",
        2467 => x"13840500",
        2468 => x"83a50500",
        2469 => x"23229100",
        2470 => x"23261100",
        2471 => x"93040500",
        2472 => x"63840500",
        2473 => x"eff01ffe",
        2474 => x"93050400",
        2475 => x"03248100",
        2476 => x"8320c100",
        2477 => x"13850400",
        2478 => x"83244100",
        2479 => x"13010101",
        2480 => x"6f004019",
        2481 => x"83a7c187",
        2482 => x"6382a716",
        2483 => x"83274502",
        2484 => x"130101fe",
        2485 => x"232c8100",
        2486 => x"232e1100",
        2487 => x"232a9100",
        2488 => x"23282101",
        2489 => x"23263101",
        2490 => x"13040500",
        2491 => x"638a0704",
        2492 => x"83a7c700",
        2493 => x"638c0702",
        2494 => x"93040000",
        2495 => x"13090008",
        2496 => x"83274402",
        2497 => x"83a7c700",
        2498 => x"b3879700",
        2499 => x"83a50700",
        2500 => x"6396050e",
        2501 => x"93844400",
        2502 => x"e39424ff",
        2503 => x"83274402",
        2504 => x"13050400",
        2505 => x"83a5c700",
        2506 => x"ef00c012",
        2507 => x"83274402",
        2508 => x"83a50700",
        2509 => x"63860500",
        2510 => x"13050400",
        2511 => x"ef008011",
        2512 => x"83254401",
        2513 => x"63860500",
        2514 => x"13050400",
        2515 => x"ef008010",
        2516 => x"83254402",
        2517 => x"63860500",
        2518 => x"13050400",
        2519 => x"ef00800f",
        2520 => x"83258403",
        2521 => x"63860500",
        2522 => x"13050400",
        2523 => x"ef00800e",
        2524 => x"8325c403",
        2525 => x"63860500",
        2526 => x"13050400",
        2527 => x"ef00800d",
        2528 => x"83250404",
        2529 => x"63860500",
        2530 => x"13050400",
        2531 => x"ef00800c",
        2532 => x"8325c405",
        2533 => x"63860500",
        2534 => x"13050400",
        2535 => x"ef00800b",
        2536 => x"83258405",
        2537 => x"63860500",
        2538 => x"13050400",
        2539 => x"ef00800a",
        2540 => x"83254403",
        2541 => x"63860500",
        2542 => x"13050400",
        2543 => x"ef008009",
        2544 => x"83278401",
        2545 => x"63860704",
        2546 => x"83278402",
        2547 => x"13050400",
        2548 => x"e7800700",
        2549 => x"83258404",
        2550 => x"638c0502",
        2551 => x"13050400",
        2552 => x"03248101",
        2553 => x"8320c101",
        2554 => x"83244101",
        2555 => x"03290101",
        2556 => x"8329c100",
        2557 => x"13010102",
        2558 => x"6ff0dfe8",
        2559 => x"83a90500",
        2560 => x"13050400",
        2561 => x"ef000005",
        2562 => x"93850900",
        2563 => x"6ff05ff0",
        2564 => x"8320c101",
        2565 => x"03248101",
        2566 => x"83244101",
        2567 => x"03290101",
        2568 => x"8329c100",
        2569 => x"13010102",
        2570 => x"67800000",
        2571 => x"67800000",
        2572 => x"93f5f50f",
        2573 => x"3306c500",
        2574 => x"6316c500",
        2575 => x"13050000",
        2576 => x"67800000",
        2577 => x"83470500",
        2578 => x"e38cb7fe",
        2579 => x"13051500",
        2580 => x"6ff09ffe",
        2581 => x"638a050e",
        2582 => x"83a7c5ff",
        2583 => x"130101fe",
        2584 => x"232c8100",
        2585 => x"232e1100",
        2586 => x"1384c5ff",
        2587 => x"63d40700",
        2588 => x"3304f400",
        2589 => x"2326a100",
        2590 => x"ef008033",
        2591 => x"83a70189",
        2592 => x"0325c100",
        2593 => x"639e0700",
        2594 => x"23220400",
        2595 => x"23a88188",
        2596 => x"03248101",
        2597 => x"8320c101",
        2598 => x"13010102",
        2599 => x"6f008031",
        2600 => x"6374f402",
        2601 => x"03260400",
        2602 => x"b306c400",
        2603 => x"639ad700",
        2604 => x"83a60700",
        2605 => x"83a74700",
        2606 => x"b386c600",
        2607 => x"2320d400",
        2608 => x"2322f400",
        2609 => x"6ff09ffc",
        2610 => x"13870700",
        2611 => x"83a74700",
        2612 => x"63840700",
        2613 => x"e37af4fe",
        2614 => x"83260700",
        2615 => x"3306d700",
        2616 => x"63188602",
        2617 => x"03260400",
        2618 => x"b386c600",
        2619 => x"2320d700",
        2620 => x"3306d700",
        2621 => x"e39ec7f8",
        2622 => x"03a60700",
        2623 => x"83a74700",
        2624 => x"b306d600",
        2625 => x"2320d700",
        2626 => x"2322f700",
        2627 => x"6ff05ff8",
        2628 => x"6378c400",
        2629 => x"9307c000",
        2630 => x"2320f500",
        2631 => x"6ff05ff7",
        2632 => x"03260400",
        2633 => x"b306c400",
        2634 => x"639ad700",
        2635 => x"83a60700",
        2636 => x"83a74700",
        2637 => x"b386c600",
        2638 => x"2320d400",
        2639 => x"2322f400",
        2640 => x"23228700",
        2641 => x"6ff0dff4",
        2642 => x"67800000",
        2643 => x"130101fe",
        2644 => x"232a9100",
        2645 => x"93843500",
        2646 => x"93f4c4ff",
        2647 => x"23282101",
        2648 => x"232e1100",
        2649 => x"232c8100",
        2650 => x"23263101",
        2651 => x"93848400",
        2652 => x"9307c000",
        2653 => x"13090500",
        2654 => x"63f0f406",
        2655 => x"9304c000",
        2656 => x"63eeb404",
        2657 => x"13050900",
        2658 => x"ef008022",
        2659 => x"03a70189",
        2660 => x"13040700",
        2661 => x"63180406",
        2662 => x"83a7c188",
        2663 => x"639a0700",
        2664 => x"93050000",
        2665 => x"13050900",
        2666 => x"ef00001c",
        2667 => x"23a6a188",
        2668 => x"93850400",
        2669 => x"13050900",
        2670 => x"ef00001b",
        2671 => x"9309f0ff",
        2672 => x"631a350b",
        2673 => x"9307c000",
        2674 => x"2320f900",
        2675 => x"13050900",
        2676 => x"ef00401e",
        2677 => x"6f000001",
        2678 => x"e3d404fa",
        2679 => x"9307c000",
        2680 => x"2320f900",
        2681 => x"13050000",
        2682 => x"8320c101",
        2683 => x"03248101",
        2684 => x"83244101",
        2685 => x"03290101",
        2686 => x"8329c100",
        2687 => x"13010102",
        2688 => x"67800000",
        2689 => x"83270400",
        2690 => x"b3879740",
        2691 => x"63ce0704",
        2692 => x"1306b000",
        2693 => x"637af600",
        2694 => x"2320f400",
        2695 => x"3304f400",
        2696 => x"23209400",
        2697 => x"6f000001",
        2698 => x"83274400",
        2699 => x"631a8702",
        2700 => x"23a8f188",
        2701 => x"13050900",
        2702 => x"ef00c017",
        2703 => x"1305b400",
        2704 => x"93074400",
        2705 => x"137585ff",
        2706 => x"3307f540",
        2707 => x"e30ef5f8",
        2708 => x"3304e400",
        2709 => x"b387a740",
        2710 => x"2320f400",
        2711 => x"6ff0dff8",
        2712 => x"2322f700",
        2713 => x"6ff01ffd",
        2714 => x"13070400",
        2715 => x"03244400",
        2716 => x"6ff05ff2",
        2717 => x"13043500",
        2718 => x"1374c4ff",
        2719 => x"e30285fa",
        2720 => x"b305a440",
        2721 => x"13050900",
        2722 => x"ef00000e",
        2723 => x"e31a35f9",
        2724 => x"6ff05ff3",
        2725 => x"130101fe",
        2726 => x"232c8100",
        2727 => x"232e1100",
        2728 => x"232a9100",
        2729 => x"23282101",
        2730 => x"23263101",
        2731 => x"23244101",
        2732 => x"13040600",
        2733 => x"63940502",
        2734 => x"03248101",
        2735 => x"8320c101",
        2736 => x"83244101",
        2737 => x"03290101",
        2738 => x"8329c100",
        2739 => x"032a8100",
        2740 => x"93050600",
        2741 => x"13010102",
        2742 => x"6ff05fe7",
        2743 => x"63180602",
        2744 => x"eff05fd7",
        2745 => x"93040000",
        2746 => x"8320c101",
        2747 => x"03248101",
        2748 => x"03290101",
        2749 => x"8329c100",
        2750 => x"032a8100",
        2751 => x"13850400",
        2752 => x"83244101",
        2753 => x"13010102",
        2754 => x"67800000",
        2755 => x"130a0500",
        2756 => x"93840500",
        2757 => x"ef00400a",
        2758 => x"13090500",
        2759 => x"63668500",
        2760 => x"93571500",
        2761 => x"e3e287fc",
        2762 => x"93050400",
        2763 => x"13050a00",
        2764 => x"eff0dfe1",
        2765 => x"93090500",
        2766 => x"e30605fa",
        2767 => x"13060400",
        2768 => x"63748900",
        2769 => x"13060900",
        2770 => x"93850400",
        2771 => x"13850900",
        2772 => x"efe08ffc",
        2773 => x"93850400",
        2774 => x"13050a00",
        2775 => x"eff09fcf",
        2776 => x"93840900",
        2777 => x"6ff05ff8",
        2778 => x"130101ff",
        2779 => x"23248100",
        2780 => x"23229100",
        2781 => x"13040500",
        2782 => x"13850500",
        2783 => x"23261100",
        2784 => x"23a40188",
        2785 => x"efe01f8a",
        2786 => x"9307f0ff",
        2787 => x"6318f500",
        2788 => x"83a78188",
        2789 => x"63840700",
        2790 => x"2320f400",
        2791 => x"8320c100",
        2792 => x"03248100",
        2793 => x"83244100",
        2794 => x"13010101",
        2795 => x"67800000",
        2796 => x"67800000",
        2797 => x"67800000",
        2798 => x"83a7c5ff",
        2799 => x"1385c7ff",
        2800 => x"63d80700",
        2801 => x"b385a500",
        2802 => x"83a70500",
        2803 => x"3305f500",
        2804 => x"67800000",
        2805 => x"10000000",
        2806 => x"00000000",
        2807 => x"037a5200",
        2808 => x"017c0101",
        2809 => x"1b0d0200",
        2810 => x"10000000",
        2811 => x"18000000",
        2812 => x"9cdaffff",
        2813 => x"78040000",
        2814 => x"00000000",
        2815 => x"10000000",
        2816 => x"00000000",
        2817 => x"037a5200",
        2818 => x"017c0101",
        2819 => x"1b0d0200",
        2820 => x"10000000",
        2821 => x"18000000",
        2822 => x"ecdeffff",
        2823 => x"30040000",
        2824 => x"00000000",
        2825 => x"10000000",
        2826 => x"00000000",
        2827 => x"037a5200",
        2828 => x"017c0101",
        2829 => x"1b0d0200",
        2830 => x"10000000",
        2831 => x"18000000",
        2832 => x"f4e2ffff",
        2833 => x"e4030000",
        2834 => x"00000000",
        2835 => x"30313233",
        2836 => x"34353637",
        2837 => x"38396162",
        2838 => x"63646566",
        2839 => x"00000000",
        2840 => x"70040000",
        2841 => x"7c040000",
        2842 => x"4c040000",
        2843 => x"64040000",
        2844 => x"58040000",
        2845 => x"8c030000",
        2846 => x"8c030000",
        2847 => x"8c030000",
        2848 => x"c0040000",
        2849 => x"8c030000",
        2850 => x"8c030000",
        2851 => x"8c030000",
        2852 => x"8c030000",
        2853 => x"8c030000",
        2854 => x"8c030000",
        2855 => x"8c030000",
        2856 => x"88040000",
        2857 => x"24050000",
        2858 => x"dc040000",
        2859 => x"dc040000",
        2860 => x"dc040000",
        2861 => x"dc040000",
        2862 => x"18050000",
        2863 => x"64050000",
        2864 => x"3c050000",
        2865 => x"dc040000",
        2866 => x"dc040000",
        2867 => x"dc040000",
        2868 => x"dc040000",
        2869 => x"dc040000",
        2870 => x"dc040000",
        2871 => x"dc040000",
        2872 => x"dc040000",
        2873 => x"dc040000",
        2874 => x"dc040000",
        2875 => x"dc040000",
        2876 => x"dc040000",
        2877 => x"dc040000",
        2878 => x"dc040000",
        2879 => x"04050000",
        2880 => x"04050000",
        2881 => x"dc040000",
        2882 => x"dc040000",
        2883 => x"dc040000",
        2884 => x"dc040000",
        2885 => x"dc040000",
        2886 => x"dc040000",
        2887 => x"dc040000",
        2888 => x"dc040000",
        2889 => x"dc040000",
        2890 => x"dc040000",
        2891 => x"dc040000",
        2892 => x"dc040000",
        2893 => x"18050000",
        2894 => x"24050000",
        2895 => x"e0050000",
        2896 => x"c8050000",
        2897 => x"dc040000",
        2898 => x"dc040000",
        2899 => x"dc040000",
        2900 => x"dc040000",
        2901 => x"dc040000",
        2902 => x"dc040000",
        2903 => x"b0050000",
        2904 => x"dc040000",
        2905 => x"dc040000",
        2906 => x"dc040000",
        2907 => x"dc040000",
        2908 => x"04050000",
        2909 => x"04050000",
        2910 => x"00010202",
        2911 => x"03030303",
        2912 => x"04040404",
        2913 => x"04040404",
        2914 => x"05050505",
        2915 => x"05050505",
        2916 => x"05050505",
        2917 => x"05050505",
        2918 => x"06060606",
        2919 => x"06060606",
        2920 => x"06060606",
        2921 => x"06060606",
        2922 => x"06060606",
        2923 => x"06060606",
        2924 => x"06060606",
        2925 => x"06060606",
        2926 => x"07070707",
        2927 => x"07070707",
        2928 => x"07070707",
        2929 => x"07070707",
        2930 => x"07070707",
        2931 => x"07070707",
        2932 => x"07070707",
        2933 => x"07070707",
        2934 => x"07070707",
        2935 => x"07070707",
        2936 => x"07070707",
        2937 => x"07070707",
        2938 => x"07070707",
        2939 => x"07070707",
        2940 => x"07070707",
        2941 => x"07070707",
        2942 => x"08080808",
        2943 => x"08080808",
        2944 => x"08080808",
        2945 => x"08080808",
        2946 => x"08080808",
        2947 => x"08080808",
        2948 => x"08080808",
        2949 => x"08080808",
        2950 => x"08080808",
        2951 => x"08080808",
        2952 => x"08080808",
        2953 => x"08080808",
        2954 => x"08080808",
        2955 => x"08080808",
        2956 => x"08080808",
        2957 => x"08080808",
        2958 => x"08080808",
        2959 => x"08080808",
        2960 => x"08080808",
        2961 => x"08080808",
        2962 => x"08080808",
        2963 => x"08080808",
        2964 => x"08080808",
        2965 => x"08080808",
        2966 => x"08080808",
        2967 => x"08080808",
        2968 => x"08080808",
        2969 => x"08080808",
        2970 => x"08080808",
        2971 => x"08080808",
        2972 => x"08080808",
        2973 => x"08080808",
        2974 => x"0d0a4542",
        2975 => x"5245414b",
        2976 => x"21206d65",
        2977 => x"7063203d",
        2978 => x"20000000",
        2979 => x"20696e73",
        2980 => x"6e203d20",
        2981 => x"00000000",
        2982 => x"0d0a0d0a",
        2983 => x"44697370",
        2984 => x"6c617969",
        2985 => x"6e672074",
        2986 => x"68652074",
        2987 => x"696d6520",
        2988 => x"70617373",
        2989 => x"65642073",
        2990 => x"696e6365",
        2991 => x"20726573",
        2992 => x"65740d0a",
        2993 => x"0d0a0000",
        2994 => x"2530356c",
        2995 => x"643a2530",
        2996 => x"366c6420",
        2997 => x"20202530",
        2998 => x"326c643a",
        2999 => x"2530326c",
        3000 => x"643a2530",
        3001 => x"326c640d",
        3002 => x"00000000",
        3003 => x"696e7465",
        3004 => x"72727570",
        3005 => x"745f6469",
        3006 => x"72656374",
        3007 => x"00000000",
        3008 => x"54485541",
        3009 => x"53205249",
        3010 => x"53432d56",
        3011 => x"20525633",
        3012 => x"32494d20",
        3013 => x"62617265",
        3014 => x"206d6574",
        3015 => x"616c2070",
        3016 => x"726f6365",
        3017 => x"73736f72",
        3018 => x"00000000",
        3019 => x"54686520",
        3020 => x"48616775",
        3021 => x"6520556e",
        3022 => x"69766572",
        3023 => x"73697479",
        3024 => x"206f6620",
        3025 => x"4170706c",
        3026 => x"69656420",
        3027 => x"53636965",
        3028 => x"6e636573",
        3029 => x"00000000",
        3030 => x"44657061",
        3031 => x"72746d65",
        3032 => x"6e74206f",
        3033 => x"6620456c",
        3034 => x"65637472",
        3035 => x"6963616c",
        3036 => x"20456e67",
        3037 => x"696e6565",
        3038 => x"72696e67",
        3039 => x"00000000",
        3040 => x"4a2e452e",
        3041 => x"4a2e206f",
        3042 => x"70206465",
        3043 => x"6e204272",
        3044 => x"6f757700",
        3045 => x"232d302b",
        3046 => x"20000000",
        3047 => x"686c4c00",
        3048 => x"65666745",
        3049 => x"46470000",
        3050 => x"30313233",
        3051 => x"34353637",
        3052 => x"38394142",
        3053 => x"43444546",
        3054 => x"00000000",
        3055 => x"30313233",
        3056 => x"34353637",
        3057 => x"38396162",
        3058 => x"63646566",
        3059 => x"00000000",
        3060 => x"50230000",
        3061 => x"70230000",
        3062 => x"1c230000",
        3063 => x"1c230000",
        3064 => x"1c230000",
        3065 => x"1c230000",
        3066 => x"70230000",
        3067 => x"1c230000",
        3068 => x"1c230000",
        3069 => x"1c230000",
        3070 => x"1c230000",
        3071 => x"88250000",
        3072 => x"04240000",
        3073 => x"f0240000",
        3074 => x"1c230000",
        3075 => x"1c230000",
        3076 => x"d0250000",
        3077 => x"1c230000",
        3078 => x"04240000",
        3079 => x"1c230000",
        3080 => x"1c230000",
        3081 => x"fc240000",
        3082 => x"18000020",
        3083 => x"ec2e0000",
        3084 => x"002f0000",
        3085 => x"2c2f0000",
        3086 => x"582f0000",
        3087 => x"802f0000",
        3088 => x"00000000",
        3089 => x"00000000",
        3090 => x"00000000",
        3091 => x"00000000",
        3092 => x"00000000",
        3093 => x"00000000",
        3094 => x"00000000",
        3095 => x"00000000",
        3096 => x"00000000",
        3097 => x"00000000",
        3098 => x"00000000",
        3099 => x"00000000",
        3100 => x"00000000",
        3101 => x"00000000",
        3102 => x"00000000",
        3103 => x"00000000",
        3104 => x"00000000",
        3105 => x"00000000",
        3106 => x"00000000",
        3107 => x"00000000",
        3108 => x"00000000",
        3109 => x"00000000",
        3110 => x"00000000",
        3111 => x"00000000",
        3112 => x"00000000",
        3113 => x"80000020",
        3114 => x"18000020",
        others => (others => '0')
    );
end package processor_common_rom;
