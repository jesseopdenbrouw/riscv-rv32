-- #################################################################################################
-- # bootloader.vhd - The bootloader ROM                                                           #
-- # ********************************************************************************************* #
-- # This file is part of the THUAS RISCV RV32 Project                                             #
-- # ********************************************************************************************* #
-- # BSD 3-Clause License                                                                          #
-- #                                                                                               #
-- # Copyright (c) 2023, Jesse op den Brouw. All rights reserved.                                  #
-- #                                                                                               #
-- # Redistribution and use in source and binary forms, with or without modification, are          #
-- # permitted provided that the following conditions are met:                                     #
-- #                                                                                               #
-- # 1. Redistributions of source code must retain the above copyright notice, this list of        #
-- #    conditions and the following disclaimer.                                                   #
-- #                                                                                               #
-- # 2. Redistributions in binary form must reproduce the above copyright notice, this list of     #
-- #    conditions and the following disclaimer in the documentation and/or other materials        #
-- #    provided with the distribution.                                                            #
-- #                                                                                               #
-- # 3. Neither the name of the copyright holder nor the names of its contributors may be used to  #
-- #    endorse or promote products derived from this software without specific prior written      #
-- #    permission.                                                                                #
-- #                                                                                               #
-- # THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND ANY EXPRESS   #
-- # OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED WARRANTIES OF               #
-- # MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE    #
-- # COPYRIGHT HOLDER OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL,     #
-- # EXEMPLARY, OR CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE #
-- # GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER CAUSED    #
-- # AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT (INCLUDING     #
-- # NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED  #
-- # OF THE POSSIBILITY OF SUCH DAMAGE.                                                            #
-- # ********************************************************************************************* #
-- # https:/github.com/jesseopdenbrouw/riscv-rv32                                                  #
-- #################################################################################################

-- This file contains the description of the bootloader ROM. The ROM
-- is placed in immutable onboard RAM blocks. A read takes two
-- clock cycles, for both instruction and data.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.processor_common.all;
use work.processor_common_rom.all;

entity bootloader is
    port (I_clk : in std_logic;
          I_areset : in std_logic;
          I_pc : in data_type;
          I_memaddress : in data_type;
          I_memsize : in memsize_type;
          I_csboot : in std_logic;
          I_stall : in std_logic;
          O_instr : out data_type;
          O_dataout : out data_type;
          --
          O_load_misaligned_error : out std_logic
         );
end entity bootloader;

architecture rtl of bootloader is

-- The bootloader ROM
signal bootrom : bootloader_type := (
           0 => x"97020000",
           1 => x"93820208",
           2 => x"73905230",
           3 => x"97010010",
           4 => x"9381417f",
           5 => x"17810010",
           6 => x"1301c1fe",
           7 => x"9387c187",
           8 => x"1387c187",
           9 => x"13060000",
          10 => x"63e4e700",
          11 => x"3386e740",
          12 => x"93050000",
          13 => x"1385c187",
          14 => x"ef000007",
          15 => x"37050020",
          16 => x"9387c187",
          17 => x"13070500",
          18 => x"13060000",
          19 => x"63e4e700",
          20 => x"3386e740",
          21 => x"b7150010",
          22 => x"9385c5f1",
          23 => x"13050500",
          24 => x"ef004002",
          25 => x"ef00d025",
          26 => x"b7050020",
          27 => x"13060000",
          28 => x"93850500",
          29 => x"13055000",
          30 => x"ef000050",
          31 => x"ef005020",
          32 => x"6f000000",
          33 => x"13030500",
          34 => x"630e0600",
          35 => x"83830500",
          36 => x"23007300",
          37 => x"1306f6ff",
          38 => x"13031300",
          39 => x"93851500",
          40 => x"e31606fe",
          41 => x"67800000",
          42 => x"13030500",
          43 => x"630a0600",
          44 => x"2300b300",
          45 => x"1306f6ff",
          46 => x"13031300",
          47 => x"e31a06fe",
          48 => x"67800000",
          49 => x"03460500",
          50 => x"83c60500",
          51 => x"13051500",
          52 => x"93851500",
          53 => x"6314d600",
          54 => x"e31606fe",
          55 => x"3305d640",
          56 => x"67800000",
          57 => x"6f000000",
          58 => x"b70700f0",
          59 => x"03a54702",
          60 => x"13754500",
          61 => x"67800000",
          62 => x"370700f0",
          63 => x"83274702",
          64 => x"93f74700",
          65 => x"e38c07fe",
          66 => x"03258702",
          67 => x"1375f50f",
          68 => x"67800000",
          69 => x"130101fd",
          70 => x"23202103",
          71 => x"37190010",
          72 => x"23248102",
          73 => x"23229102",
          74 => x"232e3101",
          75 => x"232c4101",
          76 => x"232a5101",
          77 => x"23286101",
          78 => x"23267101",
          79 => x"23248101",
          80 => x"23261102",
          81 => x"93040500",
          82 => x"13040000",
          83 => x"130949bb",
          84 => x"930a5001",
          85 => x"938bf5ff",
          86 => x"130bf007",
          87 => x"130a2000",
          88 => x"93092001",
          89 => x"371c0010",
          90 => x"eff01ff9",
          91 => x"1377f50f",
          92 => x"63c4ea0a",
          93 => x"6354ea04",
          94 => x"9307d7ff",
          95 => x"63e0f904",
          96 => x"93972700",
          97 => x"b307f900",
          98 => x"83a70700",
          99 => x"67800700",
         100 => x"630a0400",
         101 => x"1304f4ff",
         102 => x"1305f007",
         103 => x"ef004011",
         104 => x"e31a04fe",
         105 => x"eff05ff5",
         106 => x"1377f50f",
         107 => x"13040000",
         108 => x"e3d2eafc",
         109 => x"9307f007",
         110 => x"630ef70c",
         111 => x"63547405",
         112 => x"9377f50f",
         113 => x"938607fe",
         114 => x"93f6f60f",
         115 => x"1306e005",
         116 => x"e36cd6f8",
         117 => x"b3868400",
         118 => x"13050700",
         119 => x"2380f600",
         120 => x"ef00000d",
         121 => x"eff05ff1",
         122 => x"1377f50f",
         123 => x"93075001",
         124 => x"13041400",
         125 => x"e3d0e7f8",
         126 => x"9307f007",
         127 => x"6302f702",
         128 => x"e34074fd",
         129 => x"13057000",
         130 => x"ef00800a",
         131 => x"eff0dfee",
         132 => x"1377f50f",
         133 => x"e3d0eaf6",
         134 => x"e31267fb",
         135 => x"630c0406",
         136 => x"1305f007",
         137 => x"ef00c008",
         138 => x"1304f4ff",
         139 => x"6ff0dff3",
         140 => x"b3848400",
         141 => x"37150010",
         142 => x"23800400",
         143 => x"130585c3",
         144 => x"ef000009",
         145 => x"8320c102",
         146 => x"13050400",
         147 => x"03248102",
         148 => x"83244102",
         149 => x"03290102",
         150 => x"8329c101",
         151 => x"032a8101",
         152 => x"832a4101",
         153 => x"032b0101",
         154 => x"832bc100",
         155 => x"032c8100",
         156 => x"13010103",
         157 => x"67800000",
         158 => x"1305ccf0",
         159 => x"ef004005",
         160 => x"eff09fe7",
         161 => x"1377f50f",
         162 => x"13040000",
         163 => x"e3d4eaee",
         164 => x"6ff05ff2",
         165 => x"13057000",
         166 => x"ef008001",
         167 => x"6ff09ff0",
         168 => x"b70700f0",
         169 => x"23a6a702",
         170 => x"23a0b702",
         171 => x"67800000",
         172 => x"1375f50f",
         173 => x"b70700f0",
         174 => x"370700f0",
         175 => x"23a4a702",
         176 => x"83274702",
         177 => x"93f70701",
         178 => x"e38c07fe",
         179 => x"67800000",
         180 => x"630e0502",
         181 => x"130101ff",
         182 => x"23248100",
         183 => x"23261100",
         184 => x"13040500",
         185 => x"03450500",
         186 => x"630a0500",
         187 => x"13041400",
         188 => x"eff01ffc",
         189 => x"03450400",
         190 => x"e31a05fe",
         191 => x"8320c100",
         192 => x"03248100",
         193 => x"13010101",
         194 => x"67800000",
         195 => x"67800000",
         196 => x"130101fe",
         197 => x"232e1100",
         198 => x"232c8100",
         199 => x"232a9100",
         200 => x"23282101",
         201 => x"23263101",
         202 => x"23244101",
         203 => x"6358a008",
         204 => x"b7190010",
         205 => x"13090500",
         206 => x"93040000",
         207 => x"13040000",
         208 => x"938999e0",
         209 => x"130a1000",
         210 => x"6f000001",
         211 => x"3364c400",
         212 => x"93841400",
         213 => x"63029904",
         214 => x"eff01fda",
         215 => x"b387a900",
         216 => x"83c70700",
         217 => x"130605fd",
         218 => x"13144400",
         219 => x"13f74700",
         220 => x"93f64704",
         221 => x"e31c07fc",
         222 => x"93f73700",
         223 => x"e38a06fc",
         224 => x"63944701",
         225 => x"13050502",
         226 => x"130595fa",
         227 => x"93841400",
         228 => x"3364a400",
         229 => x"e31299fc",
         230 => x"8320c101",
         231 => x"13050400",
         232 => x"03248101",
         233 => x"83244101",
         234 => x"03290101",
         235 => x"8329c100",
         236 => x"032a8100",
         237 => x"13010102",
         238 => x"67800000",
         239 => x"13040000",
         240 => x"6ff09ffd",
         241 => x"83470500",
         242 => x"37160010",
         243 => x"130696e0",
         244 => x"3307f600",
         245 => x"03470700",
         246 => x"93060500",
         247 => x"13758700",
         248 => x"630e0500",
         249 => x"83c71600",
         250 => x"93861600",
         251 => x"3307f600",
         252 => x"03470700",
         253 => x"13758700",
         254 => x"e31605fe",
         255 => x"13754704",
         256 => x"630a0506",
         257 => x"13050000",
         258 => x"13031000",
         259 => x"6f000002",
         260 => x"83c71600",
         261 => x"33e5a800",
         262 => x"93861600",
         263 => x"3307f600",
         264 => x"03470700",
         265 => x"13784704",
         266 => x"63000804",
         267 => x"13784700",
         268 => x"938807fd",
         269 => x"13773700",
         270 => x"13154500",
         271 => x"e31a08fc",
         272 => x"63146700",
         273 => x"93870702",
         274 => x"938797fa",
         275 => x"33e5a700",
         276 => x"83c71600",
         277 => x"93861600",
         278 => x"3307f600",
         279 => x"03470700",
         280 => x"13784704",
         281 => x"e31408fc",
         282 => x"63840500",
         283 => x"23a0d500",
         284 => x"67800000",
         285 => x"13050000",
         286 => x"6ff01fff",
         287 => x"130101fe",
         288 => x"232e1100",
         289 => x"232c8100",
         290 => x"23220100",
         291 => x"23240100",
         292 => x"23260100",
         293 => x"63000506",
         294 => x"13040500",
         295 => x"63440504",
         296 => x"93074100",
         297 => x"9306a000",
         298 => x"93059000",
         299 => x"3377d402",
         300 => x"13850700",
         301 => x"9387f7ff",
         302 => x"13060400",
         303 => x"13070703",
         304 => x"a385e700",
         305 => x"3354d402",
         306 => x"e3e2c5fe",
         307 => x"3305d500",
         308 => x"eff01fe0",
         309 => x"8320c101",
         310 => x"03248101",
         311 => x"13010102",
         312 => x"67800000",
         313 => x"1305d002",
         314 => x"eff09fdc",
         315 => x"33048040",
         316 => x"6ff01ffb",
         317 => x"13050003",
         318 => x"eff09fdb",
         319 => x"8320c101",
         320 => x"03248101",
         321 => x"13010102",
         322 => x"67800000",
         323 => x"130101fe",
         324 => x"232e1100",
         325 => x"23220100",
         326 => x"23240100",
         327 => x"23060100",
         328 => x"9387f5ff",
         329 => x"13077000",
         330 => x"6376f700",
         331 => x"93077000",
         332 => x"93058000",
         333 => x"13074100",
         334 => x"b307f700",
         335 => x"b385b740",
         336 => x"13069003",
         337 => x"9376f500",
         338 => x"13870603",
         339 => x"6374e600",
         340 => x"13877605",
         341 => x"2380e700",
         342 => x"9387f7ff",
         343 => x"13554500",
         344 => x"e392f5fe",
         345 => x"13054100",
         346 => x"eff09fd6",
         347 => x"8320c101",
         348 => x"13010102",
         349 => x"67800000",
         350 => x"130101f8",
         351 => x"232e1106",
         352 => x"232c8106",
         353 => x"232a9106",
         354 => x"23282107",
         355 => x"23263107",
         356 => x"23244107",
         357 => x"23225107",
         358 => x"23206107",
         359 => x"232e7105",
         360 => x"232c8105",
         361 => x"232a9105",
         362 => x"2328a105",
         363 => x"2326b105",
         364 => x"732410fc",
         365 => x"63160400",
         366 => x"37e4f505",
         367 => x"13040410",
         368 => x"37c50100",
         369 => x"13050520",
         370 => x"3355a402",
         371 => x"93050000",
         372 => x"37190010",
         373 => x"370a1000",
         374 => x"b709a000",
         375 => x"93041000",
         376 => x"130afaff",
         377 => x"b70a00f0",
         378 => x"93891900",
         379 => x"1305f5ff",
         380 => x"eff01fcb",
         381 => x"37150010",
         382 => x"130505c0",
         383 => x"eff05fcd",
         384 => x"37150010",
         385 => x"130545c2",
         386 => x"eff09fcc",
         387 => x"13050400",
         388 => x"eff0dfe6",
         389 => x"130589c3",
         390 => x"eff09fcb",
         391 => x"b70700f0",
         392 => x"1307f03f",
         393 => x"23a2e700",
         394 => x"b3f74401",
         395 => x"639c0700",
         396 => x"1305a002",
         397 => x"eff0dfc7",
         398 => x"83a74a00",
         399 => x"93d71700",
         400 => x"23a2fa00",
         401 => x"eff05faa",
         402 => x"13040500",
         403 => x"631a050c",
         404 => x"93841400",
         405 => x"e39a34fd",
         406 => x"b70700f0",
         407 => x"23a20700",
         408 => x"631a0400",
         409 => x"93050000",
         410 => x"13050000",
         411 => x"eff05fc3",
         412 => x"e7000400",
         413 => x"eff05fa8",
         414 => x"93071002",
         415 => x"93040000",
         416 => x"631cf51c",
         417 => x"37140010",
         418 => x"1305c4c3",
         419 => x"eff05fc4",
         420 => x"b70900f0",
         421 => x"930a3005",
         422 => x"130ba004",
         423 => x"930b3002",
         424 => x"130a2000",
         425 => x"130ca000",
         426 => x"83a74900",
         427 => x"93c71700",
         428 => x"23a2f900",
         429 => x"eff05fa4",
         430 => x"1375f50f",
         431 => x"63185517",
         432 => x"eff09fa3",
         433 => x"937cf50f",
         434 => x"9387fcfc",
         435 => x"93f7f70f",
         436 => x"6360fa10",
         437 => x"93071003",
         438 => x"6398fc04",
         439 => x"13052000",
         440 => x"eff01fc3",
         441 => x"130dd5ff",
         442 => x"13054000",
         443 => x"eff05fc2",
         444 => x"b70d01ff",
         445 => x"930c0500",
         446 => x"330dad00",
         447 => x"938dfdff",
         448 => x"639aac05",
         449 => x"930ca000",
         450 => x"eff01f9f",
         451 => x"1375f50f",
         452 => x"e31c95ff",
         453 => x"1305c4c3",
         454 => x"eff09fbb",
         455 => x"6ff0dff8",
         456 => x"13041000",
         457 => x"6ff05ff3",
         458 => x"93072003",
         459 => x"13052000",
         460 => x"639afc00",
         461 => x"eff0dfbd",
         462 => x"130dc5ff",
         463 => x"13056000",
         464 => x"6ff0dffa",
         465 => x"eff0dfbc",
         466 => x"130db5ff",
         467 => x"13058000",
         468 => x"6ff0dff9",
         469 => x"93f5ccff",
         470 => x"13052000",
         471 => x"2326b100",
         472 => x"eff01fbb",
         473 => x"8325c100",
         474 => x"93070500",
         475 => x"b7060001",
         476 => x"3706ffff",
         477 => x"13f53c00",
         478 => x"03a70500",
         479 => x"13083000",
         480 => x"9386f6ff",
         481 => x"93081000",
         482 => x"1306f60f",
         483 => x"63064503",
         484 => x"630a0503",
         485 => x"630c1501",
         486 => x"137707f0",
         487 => x"b3e7e700",
         488 => x"23a0f500",
         489 => x"938c1c00",
         490 => x"6ff09ff5",
         491 => x"3377c700",
         492 => x"93978700",
         493 => x"6ff09ffe",
         494 => x"3377b701",
         495 => x"93970701",
         496 => x"6ff0dffd",
         497 => x"3377d700",
         498 => x"93978701",
         499 => x"6ff01ffd",
         500 => x"93879cfc",
         501 => x"93f7f70f",
         502 => x"6362fa04",
         503 => x"13052000",
         504 => x"eff01fb3",
         505 => x"93077003",
         506 => x"13058000",
         507 => x"638afc00",
         508 => x"93078003",
         509 => x"13056000",
         510 => x"6384fc00",
         511 => x"13054000",
         512 => x"eff01fb1",
         513 => x"93040500",
         514 => x"930ca000",
         515 => x"eff0df8e",
         516 => x"1375f50f",
         517 => x"e31c95ff",
         518 => x"6ff0dfef",
         519 => x"eff0df8d",
         520 => x"1375f50f",
         521 => x"e31c85ff",
         522 => x"6ff0dfee",
         523 => x"63186509",
         524 => x"1305c4c3",
         525 => x"eff0dfa9",
         526 => x"93050000",
         527 => x"13050000",
         528 => x"eff01fa6",
         529 => x"23a20900",
         530 => x"e7800400",
         531 => x"b70700f0",
         532 => x"1307a00a",
         533 => x"23a2e700",
         534 => x"130589c3",
         535 => x"b7190010",
         536 => x"eff01fa7",
         537 => x"13040000",
         538 => x"371b0010",
         539 => x"b71b0010",
         540 => x"938999e0",
         541 => x"b7170010",
         542 => x"138507c4",
         543 => x"eff05fa5",
         544 => x"93059002",
         545 => x"13054101",
         546 => x"eff0df88",
         547 => x"13054101",
         548 => x"ef00c02c",
         549 => x"b7170010",
         550 => x"130a0500",
         551 => x"938547c4",
         552 => x"13054101",
         553 => x"eff01f82",
         554 => x"631e0500",
         555 => x"37150010",
         556 => x"130585c4",
         557 => x"eff0dfa1",
         558 => x"6f004003",
         559 => x"e31c75e5",
         560 => x"6ff0dff8",
         561 => x"b7170010",
         562 => x"938547d3",
         563 => x"13054101",
         564 => x"eff04fff",
         565 => x"63100502",
         566 => x"93050000",
         567 => x"eff05f9c",
         568 => x"b70700f0",
         569 => x"23a20700",
         570 => x"e7800400",
         571 => x"e3040af8",
         572 => x"6f004018",
         573 => x"b7170010",
         574 => x"13063000",
         575 => x"938587d3",
         576 => x"13054101",
         577 => x"ef004027",
         578 => x"63100504",
         579 => x"93050000",
         580 => x"13057101",
         581 => x"eff01fab",
         582 => x"93773500",
         583 => x"13040500",
         584 => x"63940706",
         585 => x"93058000",
         586 => x"eff05fbe",
         587 => x"37150010",
         588 => x"1305c5d3",
         589 => x"eff0df99",
         590 => x"03250400",
         591 => x"93058000",
         592 => x"eff0dfbc",
         593 => x"6ff09ffa",
         594 => x"13063000",
         595 => x"93058bd5",
         596 => x"13054101",
         597 => x"ef004022",
         598 => x"631e0502",
         599 => x"93050101",
         600 => x"13057101",
         601 => x"eff01fa6",
         602 => x"93773500",
         603 => x"13040500",
         604 => x"639c0700",
         605 => x"03250101",
         606 => x"93050000",
         607 => x"eff09fa4",
         608 => x"2320a400",
         609 => x"6ff09ff6",
         610 => x"37150010",
         611 => x"130505d4",
         612 => x"6ff05ff2",
         613 => x"13063000",
         614 => x"9385cbd5",
         615 => x"13054101",
         616 => x"ef00801d",
         617 => x"83474101",
         618 => x"1307e006",
         619 => x"630c0508",
         620 => x"639ae70a",
         621 => x"93773400",
         622 => x"e39807fc",
         623 => x"130c0404",
         624 => x"b71c0010",
         625 => x"371d0010",
         626 => x"930d80ff",
         627 => x"93058000",
         628 => x"13050400",
         629 => x"eff09fb3",
         630 => x"1385ccd3",
         631 => x"eff05f8f",
         632 => x"83270400",
         633 => x"93058000",
         634 => x"130a8001",
         635 => x"13850700",
         636 => x"2326f100",
         637 => x"eff09fb1",
         638 => x"13050dd6",
         639 => x"eff05f8d",
         640 => x"b70a00ff",
         641 => x"8327c100",
         642 => x"33f55701",
         643 => x"33554501",
         644 => x"b3063501",
         645 => x"83c60600",
         646 => x"93f67609",
         647 => x"63800604",
         648 => x"130a8aff",
         649 => x"eff0df88",
         650 => x"93da8a00",
         651 => x"e31cbafd",
         652 => x"13044400",
         653 => x"130589c3",
         654 => x"eff09f89",
         655 => x"e31884f9",
         656 => x"6ff05fe3",
         657 => x"e388e7f6",
         658 => x"93050000",
         659 => x"13057101",
         660 => x"eff05f97",
         661 => x"13040500",
         662 => x"6ff0dff5",
         663 => x"1305e002",
         664 => x"6ff01ffc",
         665 => x"e3080ae0",
         666 => x"37150010",
         667 => x"130545d6",
         668 => x"eff01f86",
         669 => x"130589c3",
         670 => x"eff09f85",
         671 => x"6ff09fdf",
         672 => x"130101ff",
         673 => x"23248100",
         674 => x"23261100",
         675 => x"93070000",
         676 => x"13040500",
         677 => x"63880700",
         678 => x"93050000",
         679 => x"97000000",
         680 => x"e7000000",
         681 => x"b7170010",
         682 => x"03a587f1",
         683 => x"83278502",
         684 => x"63840700",
         685 => x"e7800700",
         686 => x"13050400",
         687 => x"eff08fe2",
         688 => x"130101ff",
         689 => x"23248100",
         690 => x"23229100",
         691 => x"37140010",
         692 => x"b7140010",
         693 => x"9387c4f1",
         694 => x"1304c4f1",
         695 => x"3304f440",
         696 => x"23202101",
         697 => x"23261100",
         698 => x"13542440",
         699 => x"9384c4f1",
         700 => x"13090000",
         701 => x"63108904",
         702 => x"b7140010",
         703 => x"37140010",
         704 => x"9387c4f1",
         705 => x"1304c4f1",
         706 => x"3304f440",
         707 => x"13542440",
         708 => x"9384c4f1",
         709 => x"13090000",
         710 => x"63188902",
         711 => x"8320c100",
         712 => x"03248100",
         713 => x"83244100",
         714 => x"03290100",
         715 => x"13010101",
         716 => x"67800000",
         717 => x"83a70400",
         718 => x"13091900",
         719 => x"93844400",
         720 => x"e7800700",
         721 => x"6ff01ffb",
         722 => x"83a70400",
         723 => x"13091900",
         724 => x"93844400",
         725 => x"e7800700",
         726 => x"6ff01ffc",
         727 => x"93070500",
         728 => x"03c70700",
         729 => x"93871700",
         730 => x"e31c07fe",
         731 => x"3385a740",
         732 => x"1305f5ff",
         733 => x"67800000",
         734 => x"630a0602",
         735 => x"1306f6ff",
         736 => x"13070000",
         737 => x"b307e500",
         738 => x"b386e500",
         739 => x"83c70700",
         740 => x"83c60600",
         741 => x"6398d700",
         742 => x"6306c700",
         743 => x"13071700",
         744 => x"e39207fe",
         745 => x"3385d740",
         746 => x"67800000",
         747 => x"13050000",
         748 => x"67800000",
         749 => x"78020010",
         750 => x"bc010010",
         751 => x"bc010010",
         752 => x"bc010010",
         753 => x"bc010010",
         754 => x"1c020010",
         755 => x"bc010010",
         756 => x"30020010",
         757 => x"bc010010",
         758 => x"bc010010",
         759 => x"30020010",
         760 => x"bc010010",
         761 => x"bc010010",
         762 => x"bc010010",
         763 => x"bc010010",
         764 => x"bc010010",
         765 => x"bc010010",
         766 => x"bc010010",
         767 => x"90010010",
         768 => x"0d0a5448",
         769 => x"55415320",
         770 => x"52495343",
         771 => x"2d562042",
         772 => x"6f6f746c",
         773 => x"6f616465",
         774 => x"72207630",
         775 => x"2e340d0a",
         776 => x"00000000",
         777 => x"436c6f63",
         778 => x"6b206672",
         779 => x"65717565",
         780 => x"6e63793a",
         781 => x"20000000",
         782 => x"0d0a0000",
         783 => x"3f0a0000",
         784 => x"3e200000",
         785 => x"68000000",
         786 => x"48656c70",
         787 => x"3a0d0a20",
         788 => x"68202020",
         789 => x"20202020",
         790 => x"20202020",
         791 => x"20202020",
         792 => x"202d2074",
         793 => x"68697320",
         794 => x"68656c70",
         795 => x"0d0a2072",
         796 => x"20202020",
         797 => x"20202020",
         798 => x"20202020",
         799 => x"20202020",
         800 => x"2d207275",
         801 => x"6e206170",
         802 => x"706c6963",
         803 => x"6174696f",
         804 => x"6e0d0a20",
         805 => x"7277203c",
         806 => x"61646472",
         807 => x"3e202020",
         808 => x"20202020",
         809 => x"202d2072",
         810 => x"65616420",
         811 => x"776f7264",
         812 => x"2066726f",
         813 => x"6d206164",
         814 => x"64720d0a",
         815 => x"20777720",
         816 => x"3c616464",
         817 => x"723e203c",
         818 => x"64617461",
         819 => x"3e202d20",
         820 => x"77726974",
         821 => x"6520776f",
         822 => x"72642064",
         823 => x"61746120",
         824 => x"61742061",
         825 => x"6464720d",
         826 => x"0a206477",
         827 => x"203c6164",
         828 => x"64723e20",
         829 => x"20202020",
         830 => x"2020202d",
         831 => x"2064756d",
         832 => x"70203136",
         833 => x"20776f72",
         834 => x"64730d0a",
         835 => x"206e2020",
         836 => x"20202020",
         837 => x"20202020",
         838 => x"20202020",
         839 => x"20202d20",
         840 => x"64756d70",
         841 => x"206e6578",
         842 => x"74203136",
         843 => x"20776f72",
         844 => x"64730000",
         845 => x"72000000",
         846 => x"72772000",
         847 => x"3a200000",
         848 => x"4e6f7420",
         849 => x"6f6e2034",
         850 => x"2d627974",
         851 => x"6520626f",
         852 => x"756e6461",
         853 => x"72792100",
         854 => x"77772000",
         855 => x"64772000",
         856 => x"20200000",
         857 => x"3f3f0000",
         858 => x"626f6f74",
         859 => x"6c6f6164",
         860 => x"65720000",
         861 => x"54485541",
         862 => x"53205249",
         863 => x"53432d56",
         864 => x"20525633",
         865 => x"32494d20",
         866 => x"62617265",
         867 => x"206d6574",
         868 => x"616c2070",
         869 => x"726f6365",
         870 => x"73736f72",
         871 => x"00000000",
         872 => x"54686520",
         873 => x"48616775",
         874 => x"6520556e",
         875 => x"69766572",
         876 => x"73697479",
         877 => x"206f6620",
         878 => x"4170706c",
         879 => x"69656420",
         880 => x"53636965",
         881 => x"6e636573",
         882 => x"00000000",
         883 => x"44657061",
         884 => x"72746d65",
         885 => x"6e74206f",
         886 => x"6620456c",
         887 => x"65637472",
         888 => x"6963616c",
         889 => x"20456e67",
         890 => x"696e6565",
         891 => x"72696e67",
         892 => x"00000000",
         893 => x"4a2e452e",
         894 => x"4a2e206f",
         895 => x"70206465",
         896 => x"6e204272",
         897 => x"6f757700",
         898 => x"00202020",
         899 => x"20202020",
         900 => x"20202828",
         901 => x"28282820",
         902 => x"20202020",
         903 => x"20202020",
         904 => x"20202020",
         905 => x"20202020",
         906 => x"20881010",
         907 => x"10101010",
         908 => x"10101010",
         909 => x"10101010",
         910 => x"10040404",
         911 => x"04040404",
         912 => x"04040410",
         913 => x"10101010",
         914 => x"10104141",
         915 => x"41414141",
         916 => x"01010101",
         917 => x"01010101",
         918 => x"01010101",
         919 => x"01010101",
         920 => x"01010101",
         921 => x"10101010",
         922 => x"10104242",
         923 => x"42424242",
         924 => x"02020202",
         925 => x"02020202",
         926 => x"02020202",
         927 => x"02020202",
         928 => x"02020202",
         929 => x"10101010",
         930 => x"20000000",
         931 => x"00000000",
         932 => x"00000000",
         933 => x"00000000",
         934 => x"00000000",
         935 => x"00000000",
         936 => x"00000000",
         937 => x"00000000",
         938 => x"00000000",
         939 => x"00000000",
         940 => x"00000000",
         941 => x"00000000",
         942 => x"00000000",
         943 => x"00000000",
         944 => x"00000000",
         945 => x"00000000",
         946 => x"00000000",
         947 => x"00000000",
         948 => x"00000000",
         949 => x"00000000",
         950 => x"00000000",
         951 => x"00000000",
         952 => x"00000000",
         953 => x"00000000",
         954 => x"00000000",
         955 => x"00000000",
         956 => x"00000000",
         957 => x"00000000",
         958 => x"00000000",
         959 => x"00000000",
         960 => x"00000000",
         961 => x"00000000",
         962 => x"00000000",
         963 => x"3c627265",
         964 => x"616b3e0d",
         965 => x"0a000000",
         966 => x"18000020",
         967 => x"680d0010",
         968 => x"740d0010",
         969 => x"a00d0010",
         970 => x"cc0d0010",
         971 => x"f40d0010",
         972 => x"00000000",
         973 => x"00000000",
         974 => x"00000000",
         975 => x"00000000",
         976 => x"00000000",
         977 => x"00000000",
         978 => x"00000000",
         979 => x"00000000",
         980 => x"00000000",
         981 => x"00000000",
         982 => x"00000000",
         983 => x"00000000",
         984 => x"00000000",
         985 => x"00000000",
         986 => x"00000000",
         987 => x"00000000",
         988 => x"00000000",
         989 => x"00000000",
         990 => x"00000000",
         991 => x"00000000",
         992 => x"00000000",
         993 => x"00000000",
         994 => x"00000000",
         995 => x"00000000",
         996 => x"00000000",
         997 => x"18000020",
         others => (others => '0')
        );

begin

    gen_bootrom: if HAVE_BOOTLOADER_ROM generate

        -- ROM, for both instructions and read-only data
        process (I_clk, I_areset, I_pc, I_memaddress, I_csboot, I_memsize, I_stall) is
        variable address_instr : integer range 0 to bootloader_size-1;
        variable address_data : integer range 0 to bootloader_size-1;
        variable instr_var : data_type;
        variable instr_recode : data_type;
        variable romdata_var : data_type;
        constant x : data_type := (others => 'X');
        begin
            -- Calculate addresses
            address_instr := to_integer(unsigned(I_pc(bootloader_size_bits-1 downto 2)));
            address_data := to_integer(unsigned(I_memaddress(bootloader_size_bits-1 downto 2)));

            -- Quartus will detect ROM table and uses onboard RAM
            -- Do not use reset, otherwise ROM will be created with ALMs
            if rising_edge(I_clk) then
                if I_stall = '0' then
                    instr_var := bootrom(address_instr);
                end if;
                romdata_var := bootrom(address_data);
            end if;
            
            -- Recode instruction
            O_instr <= instr_var(7 downto 0) & instr_var(15 downto 8) & instr_var(23 downto 16) & instr_var(31 downto 24);
            
            O_load_misaligned_error <= '0';
            
            -- By natural size, for data
            if I_csboot = '1' then
                if I_memsize = memsize_word and I_memaddress(1 downto 0) = "00" then
                    O_dataout <= romdata_var(7 downto 0) & romdata_var(15 downto 8) & romdata_var(23 downto 16) & romdata_var(31 downto 24);
                elsif I_memsize = memsize_halfword and I_memaddress(1 downto 0) = "00" then
                    O_dataout <= x(31 downto 16) & romdata_var(23 downto 16) & romdata_var(31 downto 24);
                elsif I_memsize = memsize_halfword and I_memaddress(1 downto 0) = "10" then
                    O_dataout <= x(31 downto 16) & romdata_var(7 downto 0) & romdata_var(15 downto 8);
                elsif I_memsize = memsize_byte then
                    case I_memaddress(1 downto 0) is
                        when "00" => O_dataout <= x(31 downto 8) & romdata_var(31 downto 24);
                        when "01" => O_dataout <= x(31 downto 8) & romdata_var(23 downto 16);
                        when "10" => O_dataout <= x(31 downto 8) & romdata_var(15 downto 8);
                        when "11" => O_dataout <= x(31 downto 8) & romdata_var(7 downto 0);
                        when others => O_dataout <= x; O_load_misaligned_error <= '1';
                    end case;
                else
                    -- Chip select, but not aligned
                    O_dataout <= x;
                    O_load_misaligned_error <= '1';
                end if;
            else
                -- No chip select, so no data
                O_dataout <= x;
            end if;
        end process;
    end generate;

    gen_bootrom_not: if not HAVE_BOOTLOADER_ROM generate
        O_load_misaligned_error <= '0';
        O_dataout <= (others => 'X');
        O_instr  <= (others => 'X');
    end generate;
end architecture rtl;
