-- #################################################################################################
-- # bootloader.vhd - The bootloader ROM                                                           #
-- # ********************************************************************************************* #
-- # This file is part of the THUAS RISCV RV32 Project                                             #
-- # ********************************************************************************************* #
-- # BSD 3-Clause License                                                                          #
-- #                                                                                               #
-- # Copyright (c) 2023, Jesse op den Brouw. All rights reserved.                                  #
-- #                                                                                               #
-- # Redistribution and use in source and binary forms, with or without modification, are          #
-- # permitted provided that the following conditions are met:                                     #
-- #                                                                                               #
-- # 1. Redistributions of source code must retain the above copyright notice, this list of        #
-- #    conditions and the following disclaimer.                                                   #
-- #                                                                                               #
-- # 2. Redistributions in binary form must reproduce the above copyright notice, this list of     #
-- #    conditions and the following disclaimer in the documentation and/or other materials        #
-- #    provided with the distribution.                                                            #
-- #                                                                                               #
-- # 3. Neither the name of the copyright holder nor the names of its contributors may be used to  #
-- #    endorse or promote products derived from this software without specific prior written      #
-- #    permission.                                                                                #
-- #                                                                                               #
-- # THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND ANY EXPRESS   #
-- # OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED WARRANTIES OF               #
-- # MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE    #
-- # COPYRIGHT HOLDER OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL,     #
-- # EXEMPLARY, OR CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE #
-- # GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER CAUSED    #
-- # AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT (INCLUDING     #
-- # NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED  #
-- # OF THE POSSIBILITY OF SUCH DAMAGE.                                                            #
-- # ********************************************************************************************* #
-- # https:/github.com/jesseopdenbrouw/riscv-minimal                                               #
-- #################################################################################################

-- This file contains the description of the bootloader ROM. The ROM
-- is placed in immutable onboard RAM blocks. A read takes two
-- clock cycles, for both instruction and data.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.processor_common.all;
use work.processor_common_rom.all;

entity bootloader is
    port (I_clk : in std_logic;
          I_areset : in std_logic;
          I_pc : in data_type;
          I_address : in data_type;
          I_csboot : in std_logic;
          I_size : in memsize_type;
          I_stall : in std_logic;
          O_instr : out data_type;
          O_data_out : out data_type;
          --
          O_instruction_misaligned_error : out std_logic;
          O_load_misaligned_error : out std_logic
         );
end entity bootloader;

architecture rtl of bootloader is

-- The bootloader ROM
signal bootrom : bootloader_type := (
           0 => x"97110010",
           1 => x"93810180",
           2 => x"17810010",
           3 => x"130181ff",
           4 => x"97020000",
           5 => x"93820206",
           6 => x"73905230",
           7 => x"37050020",
           8 => x"b7070020",
           9 => x"13060500",
          10 => x"93870700",
          11 => x"637af600",
          12 => x"3386c740",
          13 => x"93050000",
          14 => x"13050500",
          15 => x"ef00c047",
          16 => x"37050020",
          17 => x"b7070020",
          18 => x"13060500",
          19 => x"93870700",
          20 => x"637cf600",
          21 => x"b7150010",
          22 => x"3386c740",
          23 => x"9385c5cf",
          24 => x"13050500",
          25 => x"ef000043",
          26 => x"ef00c046",
          27 => x"6f000000",
          28 => x"6f000000",
          29 => x"b70700f0",
          30 => x"03a5c702",
          31 => x"13754500",
          32 => x"67800000",
          33 => x"370700f0",
          34 => x"8327c702",
          35 => x"93f74700",
          36 => x"e38c07fe",
          37 => x"03250702",
          38 => x"1375f50f",
          39 => x"67800000",
          40 => x"130101fd",
          41 => x"23202103",
          42 => x"37190010",
          43 => x"23248102",
          44 => x"23229102",
          45 => x"232e3101",
          46 => x"232c4101",
          47 => x"232a5101",
          48 => x"23286101",
          49 => x"23267101",
          50 => x"23248101",
          51 => x"23261102",
          52 => x"93040500",
          53 => x"13040000",
          54 => x"130909a6",
          55 => x"930a5001",
          56 => x"938bf5ff",
          57 => x"130bf007",
          58 => x"130a2000",
          59 => x"93092001",
          60 => x"371c0010",
          61 => x"eff01ff9",
          62 => x"1377f50f",
          63 => x"63c4ea0a",
          64 => x"6354ea04",
          65 => x"9307d7ff",
          66 => x"63e0f904",
          67 => x"93972700",
          68 => x"b307f900",
          69 => x"83a70700",
          70 => x"67800700",
          71 => x"630a0400",
          72 => x"1304f4ff",
          73 => x"1305f007",
          74 => x"ef004013",
          75 => x"e31a04fe",
          76 => x"eff05ff5",
          77 => x"1377f50f",
          78 => x"13040000",
          79 => x"e3d2eafc",
          80 => x"9307f007",
          81 => x"630ef70c",
          82 => x"63547405",
          83 => x"9377f50f",
          84 => x"938607fe",
          85 => x"93f6f60f",
          86 => x"1306e005",
          87 => x"e36cd6f8",
          88 => x"b3868400",
          89 => x"13050700",
          90 => x"2380f600",
          91 => x"ef00000f",
          92 => x"eff05ff1",
          93 => x"1377f50f",
          94 => x"93075001",
          95 => x"13041400",
          96 => x"e3d0e7f8",
          97 => x"9307f007",
          98 => x"6302f702",
          99 => x"e34074fd",
         100 => x"13057000",
         101 => x"ef00800c",
         102 => x"eff0dfee",
         103 => x"1377f50f",
         104 => x"e3d0eaf6",
         105 => x"e31267fb",
         106 => x"630c0406",
         107 => x"1305f007",
         108 => x"ef00c00a",
         109 => x"1304f4ff",
         110 => x"6ff0dff3",
         111 => x"b3848400",
         112 => x"37150010",
         113 => x"23800400",
         114 => x"130545ad",
         115 => x"ef00000b",
         116 => x"8320c102",
         117 => x"13050400",
         118 => x"03248102",
         119 => x"83244102",
         120 => x"03290102",
         121 => x"8329c101",
         122 => x"032a8101",
         123 => x"832a4101",
         124 => x"032b0101",
         125 => x"832bc100",
         126 => x"032c8100",
         127 => x"13010103",
         128 => x"67800000",
         129 => x"1305ccbe",
         130 => x"ef004007",
         131 => x"eff09fe7",
         132 => x"1377f50f",
         133 => x"13040000",
         134 => x"e3d4eaee",
         135 => x"6ff05ff2",
         136 => x"13057000",
         137 => x"ef008003",
         138 => x"6ff09ff0",
         139 => x"130101ff",
         140 => x"23261100",
         141 => x"ef008002",
         142 => x"8320c100",
         143 => x"13051000",
         144 => x"13010101",
         145 => x"67800000",
         146 => x"6ff0dfe3",
         147 => x"b70700f0",
         148 => x"23a2a702",
         149 => x"23a4b702",
         150 => x"67800000",
         151 => x"1375f50f",
         152 => x"b70700f0",
         153 => x"23a0a702",
         154 => x"370700f0",
         155 => x"8327c702",
         156 => x"93f70701",
         157 => x"e38c07fe",
         158 => x"67800000",
         159 => x"630e0502",
         160 => x"130101ff",
         161 => x"23248100",
         162 => x"23261100",
         163 => x"13040500",
         164 => x"03450500",
         165 => x"630a0500",
         166 => x"13041400",
         167 => x"eff01ffc",
         168 => x"03450400",
         169 => x"e31a05fe",
         170 => x"8320c100",
         171 => x"03248100",
         172 => x"13010101",
         173 => x"67800000",
         174 => x"67800000",
         175 => x"130101fe",
         176 => x"232e1100",
         177 => x"232c8100",
         178 => x"232a9100",
         179 => x"23282101",
         180 => x"23263101",
         181 => x"23244101",
         182 => x"6358a008",
         183 => x"b7190010",
         184 => x"13090500",
         185 => x"93040000",
         186 => x"13040000",
         187 => x"938999bf",
         188 => x"130a1000",
         189 => x"6f000001",
         190 => x"3364c400",
         191 => x"93841400",
         192 => x"63029904",
         193 => x"eff01fd8",
         194 => x"b387a900",
         195 => x"83c70700",
         196 => x"130605fd",
         197 => x"13144400",
         198 => x"13f74700",
         199 => x"93f64704",
         200 => x"e31c07fc",
         201 => x"93f73700",
         202 => x"e38a06fc",
         203 => x"63944701",
         204 => x"13050502",
         205 => x"130595fa",
         206 => x"93841400",
         207 => x"3364a400",
         208 => x"e31299fc",
         209 => x"8320c101",
         210 => x"13050400",
         211 => x"03248101",
         212 => x"83244101",
         213 => x"03290101",
         214 => x"8329c100",
         215 => x"032a8100",
         216 => x"13010102",
         217 => x"67800000",
         218 => x"13040000",
         219 => x"6ff09ffd",
         220 => x"83470500",
         221 => x"37160010",
         222 => x"130696bf",
         223 => x"3307f600",
         224 => x"03470700",
         225 => x"93060500",
         226 => x"13758700",
         227 => x"630e0500",
         228 => x"83c71600",
         229 => x"93861600",
         230 => x"3307f600",
         231 => x"03470700",
         232 => x"13758700",
         233 => x"e31605fe",
         234 => x"13754704",
         235 => x"630a0506",
         236 => x"13050000",
         237 => x"13031000",
         238 => x"6f000002",
         239 => x"83c71600",
         240 => x"33e5a800",
         241 => x"93861600",
         242 => x"3307f600",
         243 => x"03470700",
         244 => x"13784704",
         245 => x"63000804",
         246 => x"13784700",
         247 => x"938807fd",
         248 => x"13773700",
         249 => x"13154500",
         250 => x"e31a08fc",
         251 => x"63146700",
         252 => x"93870702",
         253 => x"938797fa",
         254 => x"33e5a700",
         255 => x"83c71600",
         256 => x"93861600",
         257 => x"3307f600",
         258 => x"03470700",
         259 => x"13784704",
         260 => x"e31408fc",
         261 => x"63840500",
         262 => x"23a0d500",
         263 => x"67800000",
         264 => x"13050000",
         265 => x"6ff01fff",
         266 => x"130101fe",
         267 => x"232e1100",
         268 => x"23220100",
         269 => x"23240100",
         270 => x"23060100",
         271 => x"9387f5ff",
         272 => x"13077000",
         273 => x"6376f700",
         274 => x"93077000",
         275 => x"93058000",
         276 => x"13074100",
         277 => x"b307f700",
         278 => x"b385b740",
         279 => x"13069003",
         280 => x"9376f500",
         281 => x"13870603",
         282 => x"6374e600",
         283 => x"13877605",
         284 => x"2380e700",
         285 => x"9387f7ff",
         286 => x"13554500",
         287 => x"e392f5fe",
         288 => x"13054100",
         289 => x"eff09fdf",
         290 => x"8320c101",
         291 => x"13010102",
         292 => x"67800000",
         293 => x"13030500",
         294 => x"630e0600",
         295 => x"83830500",
         296 => x"23007300",
         297 => x"1306f6ff",
         298 => x"13031300",
         299 => x"93851500",
         300 => x"e31606fe",
         301 => x"67800000",
         302 => x"13030500",
         303 => x"630a0600",
         304 => x"2300b300",
         305 => x"1306f6ff",
         306 => x"13031300",
         307 => x"e31a06fe",
         308 => x"67800000",
         309 => x"130101f8",
         310 => x"93050000",
         311 => x"1305101b",
         312 => x"232e1106",
         313 => x"232a9106",
         314 => x"23282107",
         315 => x"23263107",
         316 => x"23244107",
         317 => x"232c8106",
         318 => x"23225107",
         319 => x"23206107",
         320 => x"232e7105",
         321 => x"232c8105",
         322 => x"232a9105",
         323 => x"2328a105",
         324 => x"2326b105",
         325 => x"eff09fd3",
         326 => x"37150010",
         327 => x"1305c5aa",
         328 => x"eff0dfd5",
         329 => x"b70700f0",
         330 => x"1307f03f",
         331 => x"37091000",
         332 => x"b709a000",
         333 => x"23a2e700",
         334 => x"93041000",
         335 => x"1309f9ff",
         336 => x"370a00f0",
         337 => x"93891900",
         338 => x"6f004001",
         339 => x"eff09fb2",
         340 => x"13040500",
         341 => x"631a0502",
         342 => x"6382342b",
         343 => x"b3f72401",
         344 => x"93841400",
         345 => x"e39407fe",
         346 => x"1305a002",
         347 => x"eff01fcf",
         348 => x"83274a00",
         349 => x"93d71700",
         350 => x"2322fa00",
         351 => x"eff09faf",
         352 => x"13040500",
         353 => x"e30a05fc",
         354 => x"b70700f0",
         355 => x"23a20700",
         356 => x"eff05faf",
         357 => x"93071002",
         358 => x"23220100",
         359 => x"630ef526",
         360 => x"371a0010",
         361 => x"13054aad",
         362 => x"37190010",
         363 => x"eff01fcd",
         364 => x"13040000",
         365 => x"371b0010",
         366 => x"b71c0010",
         367 => x"b71a0010",
         368 => x"371c0010",
         369 => x"130999bf",
         370 => x"930980ff",
         371 => x"13058bad",
         372 => x"eff0dfca",
         373 => x"93059002",
         374 => x"13054101",
         375 => x"eff05fac",
         376 => x"13054101",
         377 => x"ef000046",
         378 => x"83474101",
         379 => x"93040500",
         380 => x"938787f9",
         381 => x"63920702",
         382 => x"83475101",
         383 => x"639e0700",
         384 => x"1385ccad",
         385 => x"eff09fc7",
         386 => x"e38204fc",
         387 => x"13054aad",
         388 => x"eff0dfc6",
         389 => x"6ff09ffb",
         390 => x"83474101",
         391 => x"9387e7f8",
         392 => x"63980702",
         393 => x"83475101",
         394 => x"63940702",
         395 => x"93050000",
         396 => x"13050000",
         397 => x"eff09fc1",
         398 => x"b70700f0",
         399 => x"23a20700",
         400 => x"83274100",
         401 => x"e7800700",
         402 => x"e38204f8",
         403 => x"6ff01ffc",
         404 => x"83474101",
         405 => x"9387e7f8",
         406 => x"639c0704",
         407 => x"83475101",
         408 => x"938797f8",
         409 => x"63960704",
         410 => x"83476101",
         411 => x"938707fe",
         412 => x"63900704",
         413 => x"93050000",
         414 => x"13057101",
         415 => x"eff05fcf",
         416 => x"93773500",
         417 => x"13040500",
         418 => x"6394070c",
         419 => x"93058000",
         420 => x"eff09fd9",
         421 => x"13858abc",
         422 => x"eff05fbe",
         423 => x"03250400",
         424 => x"93058000",
         425 => x"eff05fd8",
         426 => x"e38204f2",
         427 => x"6ff01ff6",
         428 => x"83474101",
         429 => x"938797f8",
         430 => x"63960704",
         431 => x"83475101",
         432 => x"938797f8",
         433 => x"63900704",
         434 => x"83476101",
         435 => x"938707fe",
         436 => x"639a0702",
         437 => x"93050101",
         438 => x"13057101",
         439 => x"eff05fc9",
         440 => x"93773500",
         441 => x"13040500",
         442 => x"63940706",
         443 => x"03250101",
         444 => x"93050000",
         445 => x"eff0dfc7",
         446 => x"2320a400",
         447 => x"e38804ec",
         448 => x"6ff0dff0",
         449 => x"83474101",
         450 => x"9387c7f9",
         451 => x"639c0700",
         452 => x"83475101",
         453 => x"938797f8",
         454 => x"63960700",
         455 => x"83476101",
         456 => x"938707fe",
         457 => x"03474101",
         458 => x"638e0702",
         459 => x"9307e006",
         460 => x"6306f704",
         461 => x"e38c04e8",
         462 => x"b7170010",
         463 => x"138587be",
         464 => x"eff0dfb3",
         465 => x"13054aad",
         466 => x"eff05fb3",
         467 => x"6ff01fe8",
         468 => x"b7170010",
         469 => x"1385c7bc",
         470 => x"eff05fb2",
         471 => x"e38804e6",
         472 => x"6ff0dfea",
         473 => x"9307e006",
         474 => x"630af700",
         475 => x"93050000",
         476 => x"13057101",
         477 => x"eff0dfbf",
         478 => x"13040500",
         479 => x"93773400",
         480 => x"e39807fc",
         481 => x"930b0404",
         482 => x"93058000",
         483 => x"13050400",
         484 => x"eff09fc9",
         485 => x"13858abc",
         486 => x"eff05fae",
         487 => x"83240400",
         488 => x"93058000",
         489 => x"130d8001",
         490 => x"13850400",
         491 => x"eff0dfc7",
         492 => x"13054cbe",
         493 => x"eff09fac",
         494 => x"b70d00ff",
         495 => x"33f5b401",
         496 => x"3355a501",
         497 => x"3307a900",
         498 => x"03470700",
         499 => x"13777709",
         500 => x"63140700",
         501 => x"1305e002",
         502 => x"130d8dff",
         503 => x"eff01fa8",
         504 => x"93dd8d00",
         505 => x"e31c3dfd",
         506 => x"13044400",
         507 => x"13054aad",
         508 => x"eff0dfa8",
         509 => x"e39a8bf8",
         510 => x"6ff05fdd",
         511 => x"b70400f0",
         512 => x"23a20400",
         513 => x"93050000",
         514 => x"eff05fa4",
         515 => x"23a20400",
         516 => x"e7000400",
         517 => x"6ff0dfd7",
         518 => x"b7140010",
         519 => x"138504ad",
         520 => x"eff0dfa5",
         521 => x"370400f0",
         522 => x"13093005",
         523 => x"930aa004",
         524 => x"130b3002",
         525 => x"130a2000",
         526 => x"9309a000",
         527 => x"6f004001",
         528 => x"638c5705",
         529 => x"638a6707",
         530 => x"138504ad",
         531 => x"eff01fa3",
         532 => x"83274400",
         533 => x"93c71700",
         534 => x"2322f400",
         535 => x"eff09f82",
         536 => x"9377f50f",
         537 => x"e39e27fd",
         538 => x"eff0df81",
         539 => x"937bf50f",
         540 => x"9387fbfc",
         541 => x"93f7f70f",
         542 => x"6378fa04",
         543 => x"93879bfc",
         544 => x"93f7f70f",
         545 => x"6374fa12",
         546 => x"eff0cfff",
         547 => x"9377f50f",
         548 => x"e39c37ff",
         549 => x"6ff05ffb",
         550 => x"138504ad",
         551 => x"eff01f9e",
         552 => x"93050000",
         553 => x"13050000",
         554 => x"eff05f9a",
         555 => x"83274100",
         556 => x"23220400",
         557 => x"e7800700",
         558 => x"b70700f0",
         559 => x"1307a00a",
         560 => x"23a2e700",
         561 => x"6ff0dfcd",
         562 => x"93071003",
         563 => x"638efb10",
         564 => x"93072003",
         565 => x"13052000",
         566 => x"6388fb14",
         567 => x"eff01f9e",
         568 => x"930b0500",
         569 => x"13058000",
         570 => x"eff05f9d",
         571 => x"938bbbff",
         572 => x"130d0500",
         573 => x"b38dab01",
         574 => x"63800b0a",
         575 => x"b7070001",
         576 => x"9387f7ff",
         577 => x"2324f100",
         578 => x"b707ffff",
         579 => x"b70b01ff",
         580 => x"9387f70f",
         581 => x"938bfbff",
         582 => x"930c3000",
         583 => x"130c1000",
         584 => x"2326f100",
         585 => x"6f008001",
         586 => x"630e8605",
         587 => x"b367f500",
         588 => x"23a0f500",
         589 => x"130d1d00",
         590 => x"6380ad07",
         591 => x"13052000",
         592 => x"eff0df97",
         593 => x"9375cdff",
         594 => x"13763d00",
         595 => x"83a60500",
         596 => x"93070500",
         597 => x"63004603",
         598 => x"13f506f0",
         599 => x"e31696fd",
         600 => x"03278100",
         601 => x"93978701",
         602 => x"b3f6e600",
         603 => x"b3e7d700",
         604 => x"6ff01ffc",
         605 => x"b3f67601",
         606 => x"93170501",
         607 => x"b3e7d700",
         608 => x"6ff01ffb",
         609 => x"0327c100",
         610 => x"93978700",
         611 => x"b3f6e600",
         612 => x"b3e7d700",
         613 => x"6ff0dff9",
         614 => x"930ba000",
         615 => x"eff08fee",
         616 => x"9377f50f",
         617 => x"e39c77ff",
         618 => x"6ff01fea",
         619 => x"13052000",
         620 => x"eff0df90",
         621 => x"93077003",
         622 => x"6380fb06",
         623 => x"93078003",
         624 => x"6384fb04",
         625 => x"13054000",
         626 => x"eff05f8f",
         627 => x"130d0500",
         628 => x"930ba000",
         629 => x"eff00feb",
         630 => x"9377f50f",
         631 => x"e39c77ff",
         632 => x"2322a101",
         633 => x"6ff05fe6",
         634 => x"13052000",
         635 => x"eff01f8d",
         636 => x"930b0500",
         637 => x"13054000",
         638 => x"eff05f8c",
         639 => x"938bdbff",
         640 => x"130d0500",
         641 => x"6ff01fef",
         642 => x"13056000",
         643 => x"eff01f8b",
         644 => x"130d0500",
         645 => x"6ff0dffb",
         646 => x"13058000",
         647 => x"eff01f8a",
         648 => x"130d0500",
         649 => x"6ff0dffa",
         650 => x"eff05f89",
         651 => x"930b0500",
         652 => x"13056000",
         653 => x"eff09f88",
         654 => x"938bcbff",
         655 => x"130d0500",
         656 => x"6ff05feb",
         657 => x"93070500",
         658 => x"03c70700",
         659 => x"93871700",
         660 => x"e31c07fe",
         661 => x"3385a740",
         662 => x"1305f5ff",
         663 => x"67800000",
         664 => x"04020010",
         665 => x"48010010",
         666 => x"48010010",
         667 => x"48010010",
         668 => x"48010010",
         669 => x"a8010010",
         670 => x"48010010",
         671 => x"bc010010",
         672 => x"48010010",
         673 => x"48010010",
         674 => x"bc010010",
         675 => x"48010010",
         676 => x"48010010",
         677 => x"48010010",
         678 => x"48010010",
         679 => x"48010010",
         680 => x"48010010",
         681 => x"48010010",
         682 => x"1c010010",
         683 => x"0d0a5448",
         684 => x"55415320",
         685 => x"52495343",
         686 => x"2d562042",
         687 => x"6f6f746c",
         688 => x"6f616465",
         689 => x"72207630",
         690 => x"2e320d0a",
         691 => x"00000000",
         692 => x"3f0a0000",
         693 => x"0d0a0000",
         694 => x"3e200000",
         695 => x"48656c70",
         696 => x"3a0d0a20",
         697 => x"68202020",
         698 => x"20202020",
         699 => x"20202020",
         700 => x"20202020",
         701 => x"202d2074",
         702 => x"68697320",
         703 => x"68656c70",
         704 => x"0d0a2072",
         705 => x"20202020",
         706 => x"20202020",
         707 => x"20202020",
         708 => x"20202020",
         709 => x"2d207275",
         710 => x"6e206170",
         711 => x"706c6963",
         712 => x"6174696f",
         713 => x"6e0d0a20",
         714 => x"7277203c",
         715 => x"61646472",
         716 => x"3e202020",
         717 => x"20202020",
         718 => x"202d2072",
         719 => x"65616420",
         720 => x"776f7264",
         721 => x"2066726f",
         722 => x"6d206164",
         723 => x"64720d0a",
         724 => x"20777720",
         725 => x"3c616464",
         726 => x"723e203c",
         727 => x"64617461",
         728 => x"3e202d20",
         729 => x"77726974",
         730 => x"6520776f",
         731 => x"72642064",
         732 => x"61746120",
         733 => x"61742061",
         734 => x"6464720d",
         735 => x"0a206477",
         736 => x"203c6164",
         737 => x"64723e20",
         738 => x"20202020",
         739 => x"2020202d",
         740 => x"2064756d",
         741 => x"70203136",
         742 => x"20776f72",
         743 => x"64730d0a",
         744 => x"206e2020",
         745 => x"20202020",
         746 => x"20202020",
         747 => x"20202020",
         748 => x"20202d20",
         749 => x"64756d70",
         750 => x"206e6578",
         751 => x"74203136",
         752 => x"20776f72",
         753 => x"64730000",
         754 => x"3a200000",
         755 => x"4e6f7420",
         756 => x"6f6e2034",
         757 => x"2d627974",
         758 => x"6520626f",
         759 => x"756e6461",
         760 => x"72792100",
         761 => x"20200000",
         762 => x"3f3f0000",
         763 => x"3c627265",
         764 => x"616b3e0d",
         765 => x"0a000000",
         766 => x"00202020",
         767 => x"20202020",
         768 => x"20202828",
         769 => x"28282820",
         770 => x"20202020",
         771 => x"20202020",
         772 => x"20202020",
         773 => x"20202020",
         774 => x"20881010",
         775 => x"10101010",
         776 => x"10101010",
         777 => x"10101010",
         778 => x"10040404",
         779 => x"04040404",
         780 => x"04040410",
         781 => x"10101010",
         782 => x"10104141",
         783 => x"41414141",
         784 => x"01010101",
         785 => x"01010101",
         786 => x"01010101",
         787 => x"01010101",
         788 => x"01010101",
         789 => x"10101010",
         790 => x"10104242",
         791 => x"42424242",
         792 => x"02020202",
         793 => x"02020202",
         794 => x"02020202",
         795 => x"02020202",
         796 => x"02020202",
         797 => x"10101010",
         798 => x"20000000",
         799 => x"00000000",
         800 => x"00000000",
         801 => x"00000000",
         802 => x"00000000",
         803 => x"00000000",
         804 => x"00000000",
         805 => x"00000000",
         806 => x"00000000",
         807 => x"00000000",
         808 => x"00000000",
         809 => x"00000000",
         810 => x"00000000",
         811 => x"00000000",
         812 => x"00000000",
         813 => x"00000000",
         814 => x"00000000",
         815 => x"00000000",
         816 => x"00000000",
         817 => x"00000000",
         818 => x"00000000",
         819 => x"00000000",
         820 => x"00000000",
         821 => x"00000000",
         822 => x"00000000",
         823 => x"00000000",
         824 => x"00000000",
         825 => x"00000000",
         826 => x"00000000",
         827 => x"00000000",
         828 => x"00000000",
         829 => x"00000000",
         830 => x"00000000",
         others => (others => '0')
        );

begin

    gen_bootrom: if HAVE_BOOTLOADER_ROM generate
        O_instruction_misaligned_error <= '0' when I_pc(1 downto 0) = "00" else '1';        

        -- ROM, for both instructions and read-only data
        process (I_clk, I_areset, I_pc, I_address, I_csboot, I_size, I_stall) is
        variable address_instr : integer range 0 to bootloader_size-1;
        variable address_data : integer range 0 to bootloader_size-1;
        variable instr_var : data_type;
        variable instr_recode : data_type;
        variable romdata_var : data_type;
        constant x : data_type := (others => 'X');
        begin
            -- Calculate addresses
            address_instr := to_integer(unsigned(I_pc(bootloader_size_bits-1 downto 2)));
            address_data := to_integer(unsigned(I_address(bootloader_size_bits-1 downto 2)));

            -- Quartus will detect ROM table and uses onboard RAM
            -- Do not use reset, otherwise ROM will be created with ALMs
            if rising_edge(I_clk) then
                if I_stall = '0' then
                    instr_var := bootrom(address_instr);
                end if;
                romdata_var := bootrom(address_data);
            end if;
            
            -- Recode instruction
            O_instr <= instr_var(7 downto 0) & instr_var(15 downto 8) & instr_var(23 downto 16) & instr_var(31 downto 24);
            
            O_load_misaligned_error <= '0';
            
            -- By natural size, for data
            if I_csboot = '1' then
                if I_size = memsize_word and I_address(1 downto 0) = "00" then
                    O_data_out <= romdata_var(7 downto 0) & romdata_var(15 downto 8) & romdata_var(23 downto 16) & romdata_var(31 downto 24);
                elsif I_size = memsize_halfword and I_address(1 downto 0) = "00" then
                    O_data_out <= x(31 downto 16) & romdata_var(23 downto 16) & romdata_var(31 downto 24);
                elsif I_size = memsize_halfword and I_address(1 downto 0) = "10" then
                    O_data_out <= x(31 downto 16) & romdata_var(7 downto 0) & romdata_var(15 downto 8);
                elsif I_size = memsize_byte then
                    case I_address(1 downto 0) is
                        when "00" => O_data_out <= x(31 downto 8) & romdata_var(31 downto 24);
                        when "01" => O_data_out <= x(31 downto 8) & romdata_var(23 downto 16);
                        when "10" => O_data_out <= x(31 downto 8) & romdata_var(15 downto 8);
                        when "11" => O_data_out <= x(31 downto 8) & romdata_var(7 downto 0);
                        when others => O_data_out <= x; O_load_misaligned_error <= '1';
                    end case;
                else
                    -- Chip select, but not aligned
                    O_data_out <= x;
                    O_load_misaligned_error <= '1';
                end if;
            else
                -- No chip select, so no data
                O_data_out <= x;
            end if;
        end process;
    end generate;

    gen_bootrom_not: if not HAVE_BOOTLOADER_ROM generate
        O_instruction_misaligned_error <= '0';
        O_load_misaligned_error <= '0';
        O_data_out <= (others => 'X');
        O_instr  <= (others => 'X');
    end generate;
end architecture rtl;
