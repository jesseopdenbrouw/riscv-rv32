-- #################################################################################################
-- # bootloader.vhd - The bootloader ROM                                                           #
-- # ********************************************************************************************* #
-- # This file is part of the THUAS RISCV RV32 Project                                             #
-- # ********************************************************************************************* #
-- # BSD 3-Clause License                                                                          #
-- #                                                                                               #
-- # Copyright (c) 2023, Jesse op den Brouw. All rights reserved.                                  #
-- #                                                                                               #
-- # Redistribution and use in source and binary forms, with or without modification, are          #
-- # permitted provided that the following conditions are met:                                     #
-- #                                                                                               #
-- # 1. Redistributions of source code must retain the above copyright notice, this list of        #
-- #    conditions and the following disclaimer.                                                   #
-- #                                                                                               #
-- # 2. Redistributions in binary form must reproduce the above copyright notice, this list of     #
-- #    conditions and the following disclaimer in the documentation and/or other materials        #
-- #    provided with the distribution.                                                            #
-- #                                                                                               #
-- # 3. Neither the name of the copyright holder nor the names of its contributors may be used to  #
-- #    endorse or promote products derived from this software without specific prior written      #
-- #    permission.                                                                                #
-- #                                                                                               #
-- # THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND ANY EXPRESS   #
-- # OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED WARRANTIES OF               #
-- # MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE    #
-- # COPYRIGHT HOLDER OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL,     #
-- # EXEMPLARY, OR CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE #
-- # GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER CAUSED    #
-- # AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT (INCLUDING     #
-- # NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED  #
-- # OF THE POSSIBILITY OF SUCH DAMAGE.                                                            #
-- # ********************************************************************************************* #
-- # https:/github.com/jesseopdenbrouw/riscv-minimal                                               #
-- #################################################################################################

-- This file contains the description of the bootloader ROM. The ROM
-- is placed in immutable onboard RAM blocks. A read takes two
-- clock cycles, for both instruction and data.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.processor_common.all;
use work.processor_common_rom.all;

entity bootloader is
    port (I_clk : in std_logic;
          I_areset : in std_logic;
          I_pc : in data_type;
          I_memaddress : in data_type;
          I_memsize : in memsize_type;
          I_csboot : in std_logic;
          I_stall : in std_logic;
          O_instr : out data_type;
          O_dataout : out data_type;
          --
          O_instruction_misaligned_error : out std_logic;
          O_load_misaligned_error : out std_logic
         );
end entity bootloader;

architecture rtl of bootloader is

-- The bootloader ROM
signal bootrom : bootloader_type := (
           0 => x"97020000",
           1 => x"93820208",
           2 => x"73905230",
           3 => x"97010010",
           4 => x"9381417f",
           5 => x"17810010",
           6 => x"1301c1fe",
           7 => x"9387c187",
           8 => x"1387c187",
           9 => x"13060000",
          10 => x"63e4e700",
          11 => x"3386e740",
          12 => x"93050000",
          13 => x"1385c187",
          14 => x"ef000047",
          15 => x"37050020",
          16 => x"9387c187",
          17 => x"13070500",
          18 => x"13060000",
          19 => x"63e4e700",
          20 => x"3386e740",
          21 => x"b7150010",
          22 => x"9385c5e3",
          23 => x"13050500",
          24 => x"ef004042",
          25 => x"ef005019",
          26 => x"b7050020",
          27 => x"13060000",
          28 => x"93850500",
          29 => x"13055000",
          30 => x"ef000047",
          31 => x"ef00d013",
          32 => x"6f000000",
          33 => x"b70700f0",
          34 => x"03a54702",
          35 => x"13754500",
          36 => x"67800000",
          37 => x"370700f0",
          38 => x"83274702",
          39 => x"93f74700",
          40 => x"e38c07fe",
          41 => x"03258702",
          42 => x"1375f50f",
          43 => x"67800000",
          44 => x"130101fd",
          45 => x"23202103",
          46 => x"37190010",
          47 => x"23248102",
          48 => x"23229102",
          49 => x"232e3101",
          50 => x"232c4101",
          51 => x"232a5101",
          52 => x"23286101",
          53 => x"23267101",
          54 => x"23248101",
          55 => x"23261102",
          56 => x"93040500",
          57 => x"13040000",
          58 => x"1309c9ae",
          59 => x"930a5001",
          60 => x"938bf5ff",
          61 => x"130bf007",
          62 => x"130a2000",
          63 => x"93092001",
          64 => x"371c0010",
          65 => x"eff01ff9",
          66 => x"1377f50f",
          67 => x"63c4ea0a",
          68 => x"6354ea04",
          69 => x"9307d7ff",
          70 => x"63e0f904",
          71 => x"93972700",
          72 => x"b307f900",
          73 => x"83a70700",
          74 => x"67800700",
          75 => x"630a0400",
          76 => x"1304f4ff",
          77 => x"1305f007",
          78 => x"ef004011",
          79 => x"e31a04fe",
          80 => x"eff05ff5",
          81 => x"1377f50f",
          82 => x"13040000",
          83 => x"e3d2eafc",
          84 => x"9307f007",
          85 => x"630ef70c",
          86 => x"63547405",
          87 => x"9377f50f",
          88 => x"938607fe",
          89 => x"93f6f60f",
          90 => x"1306e005",
          91 => x"e36cd6f8",
          92 => x"b3868400",
          93 => x"13050700",
          94 => x"2380f600",
          95 => x"ef00000d",
          96 => x"eff05ff1",
          97 => x"1377f50f",
          98 => x"93075001",
          99 => x"13041400",
         100 => x"e3d0e7f8",
         101 => x"9307f007",
         102 => x"6302f702",
         103 => x"e34074fd",
         104 => x"13057000",
         105 => x"ef00800a",
         106 => x"eff0dfee",
         107 => x"1377f50f",
         108 => x"e3d0eaf6",
         109 => x"e31267fb",
         110 => x"630c0406",
         111 => x"1305f007",
         112 => x"ef00c008",
         113 => x"1304f4ff",
         114 => x"6ff0dff3",
         115 => x"b3848400",
         116 => x"37150010",
         117 => x"23800400",
         118 => x"130585b5",
         119 => x"ef000009",
         120 => x"8320c102",
         121 => x"13050400",
         122 => x"03248102",
         123 => x"83244102",
         124 => x"03290102",
         125 => x"8329c101",
         126 => x"032a8101",
         127 => x"832a4101",
         128 => x"032b0101",
         129 => x"832bc100",
         130 => x"032c8100",
         131 => x"13010103",
         132 => x"67800000",
         133 => x"13058cd2",
         134 => x"ef004005",
         135 => x"eff09fe7",
         136 => x"1377f50f",
         137 => x"13040000",
         138 => x"e3d4eaee",
         139 => x"6ff05ff2",
         140 => x"13057000",
         141 => x"ef008001",
         142 => x"6ff09ff0",
         143 => x"b70700f0",
         144 => x"23a6a702",
         145 => x"23a0b702",
         146 => x"67800000",
         147 => x"1375f50f",
         148 => x"b70700f0",
         149 => x"370700f0",
         150 => x"23a4a702",
         151 => x"83274702",
         152 => x"93f70701",
         153 => x"e38c07fe",
         154 => x"67800000",
         155 => x"630e0502",
         156 => x"130101ff",
         157 => x"23248100",
         158 => x"23261100",
         159 => x"13040500",
         160 => x"03450500",
         161 => x"630a0500",
         162 => x"13041400",
         163 => x"eff01ffc",
         164 => x"03450400",
         165 => x"e31a05fe",
         166 => x"8320c100",
         167 => x"03248100",
         168 => x"13010101",
         169 => x"67800000",
         170 => x"67800000",
         171 => x"130101fe",
         172 => x"232e1100",
         173 => x"232c8100",
         174 => x"232a9100",
         175 => x"23282101",
         176 => x"23263101",
         177 => x"23244101",
         178 => x"6358a008",
         179 => x"b7190010",
         180 => x"13090500",
         181 => x"93040000",
         182 => x"13040000",
         183 => x"938959d3",
         184 => x"130a1000",
         185 => x"6f000001",
         186 => x"3364c400",
         187 => x"93841400",
         188 => x"63029904",
         189 => x"eff01fda",
         190 => x"b387a900",
         191 => x"83c70700",
         192 => x"130605fd",
         193 => x"13144400",
         194 => x"13f74700",
         195 => x"93f64704",
         196 => x"e31c07fc",
         197 => x"93f73700",
         198 => x"e38a06fc",
         199 => x"63944701",
         200 => x"13050502",
         201 => x"130595fa",
         202 => x"93841400",
         203 => x"3364a400",
         204 => x"e31299fc",
         205 => x"8320c101",
         206 => x"13050400",
         207 => x"03248101",
         208 => x"83244101",
         209 => x"03290101",
         210 => x"8329c100",
         211 => x"032a8100",
         212 => x"13010102",
         213 => x"67800000",
         214 => x"13040000",
         215 => x"6ff09ffd",
         216 => x"83470500",
         217 => x"37160010",
         218 => x"130656d3",
         219 => x"3307f600",
         220 => x"03470700",
         221 => x"93060500",
         222 => x"13758700",
         223 => x"630e0500",
         224 => x"83c71600",
         225 => x"93861600",
         226 => x"3307f600",
         227 => x"03470700",
         228 => x"13758700",
         229 => x"e31605fe",
         230 => x"13754704",
         231 => x"630a0506",
         232 => x"13050000",
         233 => x"13031000",
         234 => x"6f000002",
         235 => x"83c71600",
         236 => x"33e5a800",
         237 => x"93861600",
         238 => x"3307f600",
         239 => x"03470700",
         240 => x"13784704",
         241 => x"63000804",
         242 => x"13784700",
         243 => x"938807fd",
         244 => x"13773700",
         245 => x"13154500",
         246 => x"e31a08fc",
         247 => x"63146700",
         248 => x"93870702",
         249 => x"938797fa",
         250 => x"33e5a700",
         251 => x"83c71600",
         252 => x"93861600",
         253 => x"3307f600",
         254 => x"03470700",
         255 => x"13784704",
         256 => x"e31408fc",
         257 => x"63840500",
         258 => x"23a0d500",
         259 => x"67800000",
         260 => x"13050000",
         261 => x"6ff01fff",
         262 => x"130101fe",
         263 => x"232e1100",
         264 => x"23220100",
         265 => x"23240100",
         266 => x"23060100",
         267 => x"9387f5ff",
         268 => x"13077000",
         269 => x"6376f700",
         270 => x"93077000",
         271 => x"93058000",
         272 => x"13074100",
         273 => x"b307f700",
         274 => x"b385b740",
         275 => x"13069003",
         276 => x"9376f500",
         277 => x"13870603",
         278 => x"6374e600",
         279 => x"13877605",
         280 => x"2380e700",
         281 => x"9387f7ff",
         282 => x"13554500",
         283 => x"e392f5fe",
         284 => x"13054100",
         285 => x"eff09fdf",
         286 => x"8320c101",
         287 => x"13010102",
         288 => x"67800000",
         289 => x"13030500",
         290 => x"630e0600",
         291 => x"83830500",
         292 => x"23007300",
         293 => x"1306f6ff",
         294 => x"13031300",
         295 => x"93851500",
         296 => x"e31606fe",
         297 => x"67800000",
         298 => x"13030500",
         299 => x"630a0600",
         300 => x"2300b300",
         301 => x"1306f6ff",
         302 => x"13031300",
         303 => x"e31a06fe",
         304 => x"67800000",
         305 => x"03460500",
         306 => x"83c60500",
         307 => x"13051500",
         308 => x"93851500",
         309 => x"6314d600",
         310 => x"e31606fe",
         311 => x"3305d640",
         312 => x"67800000",
         313 => x"6f000000",
         314 => x"130101f8",
         315 => x"93050000",
         316 => x"1305101b",
         317 => x"232e1106",
         318 => x"232a9106",
         319 => x"23282107",
         320 => x"23263107",
         321 => x"23244107",
         322 => x"232c8106",
         323 => x"23225107",
         324 => x"23206107",
         325 => x"232e7105",
         326 => x"232c8105",
         327 => x"232a9105",
         328 => x"2328a105",
         329 => x"2326b105",
         330 => x"eff05fd1",
         331 => x"37150010",
         332 => x"130585b3",
         333 => x"eff09fd3",
         334 => x"b70700f0",
         335 => x"1307f03f",
         336 => x"b7091000",
         337 => x"3709a000",
         338 => x"23a2e700",
         339 => x"93041000",
         340 => x"9389f9ff",
         341 => x"370a00f0",
         342 => x"13091900",
         343 => x"b3f73401",
         344 => x"639c0700",
         345 => x"1305a002",
         346 => x"eff05fce",
         347 => x"83274a00",
         348 => x"93d71700",
         349 => x"2322fa00",
         350 => x"eff0dfb0",
         351 => x"13040500",
         352 => x"631e050c",
         353 => x"93841400",
         354 => x"e39a24fd",
         355 => x"b70700f0",
         356 => x"23a20700",
         357 => x"631a0400",
         358 => x"93050000",
         359 => x"13050000",
         360 => x"eff0dfc9",
         361 => x"e7000400",
         362 => x"eff0dfae",
         363 => x"93071002",
         364 => x"93040000",
         365 => x"631cf51c",
         366 => x"37140010",
         367 => x"1305c4b5",
         368 => x"eff0dfca",
         369 => x"370900f0",
         370 => x"130a3005",
         371 => x"930aa004",
         372 => x"130b3002",
         373 => x"93092000",
         374 => x"930ba000",
         375 => x"83274900",
         376 => x"93c71700",
         377 => x"2322f900",
         378 => x"eff0dfaa",
         379 => x"1375f50f",
         380 => x"63184517",
         381 => x"eff01faa",
         382 => x"137cf50f",
         383 => x"9307fcfc",
         384 => x"93f7f70f",
         385 => x"63e0f910",
         386 => x"93071003",
         387 => x"631cfc04",
         388 => x"13052000",
         389 => x"eff09fc9",
         390 => x"930cd5ff",
         391 => x"13054000",
         392 => x"eff0dfc8",
         393 => x"370d01ff",
         394 => x"b70d0001",
         395 => x"130c0500",
         396 => x"b38cac00",
         397 => x"130dfdff",
         398 => x"938dfdff",
         399 => x"631a9c05",
         400 => x"130ca000",
         401 => x"eff01fa5",
         402 => x"1375f50f",
         403 => x"e31c85ff",
         404 => x"1305c4b5",
         405 => x"eff09fc1",
         406 => x"6ff05ff8",
         407 => x"13041000",
         408 => x"6ff0dff2",
         409 => x"93072003",
         410 => x"13052000",
         411 => x"631afc00",
         412 => x"eff0dfc3",
         413 => x"930cc5ff",
         414 => x"13056000",
         415 => x"6ff05ffa",
         416 => x"eff0dfc2",
         417 => x"930cb5ff",
         418 => x"13058000",
         419 => x"6ff05ff9",
         420 => x"1376ccff",
         421 => x"13052000",
         422 => x"2326c100",
         423 => x"eff01fc1",
         424 => x"0326c100",
         425 => x"93070500",
         426 => x"b706ffff",
         427 => x"13753c00",
         428 => x"03270600",
         429 => x"93053000",
         430 => x"13081000",
         431 => x"9386f60f",
         432 => x"63063503",
         433 => x"630ab502",
         434 => x"630c0501",
         435 => x"137707f0",
         436 => x"b3e7e700",
         437 => x"2320f600",
         438 => x"130c1c00",
         439 => x"6ff01ff6",
         440 => x"3377d700",
         441 => x"93978700",
         442 => x"6ff09ffe",
         443 => x"3377a701",
         444 => x"93970701",
         445 => x"6ff0dffd",
         446 => x"3377b701",
         447 => x"93978701",
         448 => x"6ff01ffd",
         449 => x"93079cfc",
         450 => x"93f7f70f",
         451 => x"63e2f904",
         452 => x"13052000",
         453 => x"eff09fb9",
         454 => x"93077003",
         455 => x"13058000",
         456 => x"630afc00",
         457 => x"93078003",
         458 => x"13056000",
         459 => x"6304fc00",
         460 => x"13054000",
         461 => x"eff09fb7",
         462 => x"93040500",
         463 => x"130ca000",
         464 => x"eff05f95",
         465 => x"1375f50f",
         466 => x"e31c85ff",
         467 => x"6ff05ff0",
         468 => x"eff05f94",
         469 => x"1375f50f",
         470 => x"e31c75ff",
         471 => x"6ff05fef",
         472 => x"631a5509",
         473 => x"1305c4b5",
         474 => x"eff05fb0",
         475 => x"93050000",
         476 => x"13050000",
         477 => x"eff09fac",
         478 => x"23220900",
         479 => x"e7800400",
         480 => x"b70700f0",
         481 => x"1307a00a",
         482 => x"23a2e700",
         483 => x"37190010",
         484 => x"130589b5",
         485 => x"b7190010",
         486 => x"eff05fad",
         487 => x"13040000",
         488 => x"371b0010",
         489 => x"b71b0010",
         490 => x"938959d3",
         491 => x"b7170010",
         492 => x"138507b6",
         493 => x"eff09fab",
         494 => x"93059002",
         495 => x"13054101",
         496 => x"eff01f8f",
         497 => x"13054101",
         498 => x"ef00c02c",
         499 => x"b7170010",
         500 => x"130a0500",
         501 => x"938547b6",
         502 => x"13054101",
         503 => x"eff09fce",
         504 => x"631e0500",
         505 => x"37150010",
         506 => x"130585b6",
         507 => x"eff01fa8",
         508 => x"6f004003",
         509 => x"e31e65e5",
         510 => x"6ff09ff8",
         511 => x"b7170010",
         512 => x"938547c5",
         513 => x"13054101",
         514 => x"eff0dfcb",
         515 => x"63100502",
         516 => x"93050000",
         517 => x"eff09fa2",
         518 => x"b70700f0",
         519 => x"23a20700",
         520 => x"e7800400",
         521 => x"e3040af8",
         522 => x"6f004018",
         523 => x"b7170010",
         524 => x"13063000",
         525 => x"938587c5",
         526 => x"13054101",
         527 => x"ef004027",
         528 => x"63100504",
         529 => x"93050000",
         530 => x"13057101",
         531 => x"eff05fb1",
         532 => x"93773500",
         533 => x"13040500",
         534 => x"63940706",
         535 => x"93058000",
         536 => x"eff09fbb",
         537 => x"37150010",
         538 => x"1305c5c5",
         539 => x"eff01fa0",
         540 => x"03250400",
         541 => x"93058000",
         542 => x"eff01fba",
         543 => x"6ff09ffa",
         544 => x"13063000",
         545 => x"93058bc7",
         546 => x"13054101",
         547 => x"ef004022",
         548 => x"631e0502",
         549 => x"93050101",
         550 => x"13057101",
         551 => x"eff05fac",
         552 => x"93773500",
         553 => x"13040500",
         554 => x"639c0700",
         555 => x"03250101",
         556 => x"93050000",
         557 => x"eff0dfaa",
         558 => x"2320a400",
         559 => x"6ff09ff6",
         560 => x"37150010",
         561 => x"130505c6",
         562 => x"6ff05ff2",
         563 => x"13063000",
         564 => x"9385cbc7",
         565 => x"13054101",
         566 => x"ef00801d",
         567 => x"83474101",
         568 => x"1307e006",
         569 => x"630c0508",
         570 => x"639ae70a",
         571 => x"93773400",
         572 => x"e39807fc",
         573 => x"130c0404",
         574 => x"b71c0010",
         575 => x"371d0010",
         576 => x"930d80ff",
         577 => x"93058000",
         578 => x"13050400",
         579 => x"eff0dfb0",
         580 => x"1385ccc5",
         581 => x"eff09f95",
         582 => x"83270400",
         583 => x"93058000",
         584 => x"130a8001",
         585 => x"13850700",
         586 => x"2326f100",
         587 => x"eff0dfae",
         588 => x"13050dc8",
         589 => x"eff09f93",
         590 => x"b70a00ff",
         591 => x"8327c100",
         592 => x"33f55701",
         593 => x"33554501",
         594 => x"b3063501",
         595 => x"83c60600",
         596 => x"93f67609",
         597 => x"63800604",
         598 => x"130a8aff",
         599 => x"eff01f8f",
         600 => x"93da8a00",
         601 => x"e31cbafd",
         602 => x"13044400",
         603 => x"130589b5",
         604 => x"eff0df8f",
         605 => x"e31884f9",
         606 => x"6ff05fe3",
         607 => x"e388e7f6",
         608 => x"93050000",
         609 => x"13057101",
         610 => x"eff09f9d",
         611 => x"13040500",
         612 => x"6ff0dff5",
         613 => x"1305e002",
         614 => x"6ff01ffc",
         615 => x"e3080ae0",
         616 => x"37150010",
         617 => x"130545c8",
         618 => x"eff05f8c",
         619 => x"130589b5",
         620 => x"eff0df8b",
         621 => x"6ff09fdf",
         622 => x"130101ff",
         623 => x"23248100",
         624 => x"23261100",
         625 => x"93070000",
         626 => x"13040500",
         627 => x"63880700",
         628 => x"93050000",
         629 => x"97000000",
         630 => x"e7000000",
         631 => x"b7170010",
         632 => x"03a587e3",
         633 => x"83278502",
         634 => x"63840700",
         635 => x"e7800700",
         636 => x"13050400",
         637 => x"eff01faf",
         638 => x"130101ff",
         639 => x"23248100",
         640 => x"23229100",
         641 => x"37140010",
         642 => x"b7140010",
         643 => x"9387c4e3",
         644 => x"1304c4e3",
         645 => x"3304f440",
         646 => x"23202101",
         647 => x"23261100",
         648 => x"13542440",
         649 => x"9384c4e3",
         650 => x"13090000",
         651 => x"63108904",
         652 => x"b7140010",
         653 => x"37140010",
         654 => x"9387c4e3",
         655 => x"1304c4e3",
         656 => x"3304f440",
         657 => x"13542440",
         658 => x"9384c4e3",
         659 => x"13090000",
         660 => x"63188902",
         661 => x"8320c100",
         662 => x"03248100",
         663 => x"83244100",
         664 => x"03290100",
         665 => x"13010101",
         666 => x"67800000",
         667 => x"83a70400",
         668 => x"13091900",
         669 => x"93844400",
         670 => x"e7800700",
         671 => x"6ff01ffb",
         672 => x"83a70400",
         673 => x"13091900",
         674 => x"93844400",
         675 => x"e7800700",
         676 => x"6ff01ffc",
         677 => x"93070500",
         678 => x"03c70700",
         679 => x"93871700",
         680 => x"e31c07fe",
         681 => x"3385a740",
         682 => x"1305f5ff",
         683 => x"67800000",
         684 => x"630a0602",
         685 => x"1306f6ff",
         686 => x"13070000",
         687 => x"b307e500",
         688 => x"b386e500",
         689 => x"83c70700",
         690 => x"83c60600",
         691 => x"6398d700",
         692 => x"6306c700",
         693 => x"13071700",
         694 => x"e39207fe",
         695 => x"3385d740",
         696 => x"67800000",
         697 => x"13050000",
         698 => x"67800000",
         699 => x"14020010",
         700 => x"58010010",
         701 => x"58010010",
         702 => x"58010010",
         703 => x"58010010",
         704 => x"b8010010",
         705 => x"58010010",
         706 => x"cc010010",
         707 => x"58010010",
         708 => x"58010010",
         709 => x"cc010010",
         710 => x"58010010",
         711 => x"58010010",
         712 => x"58010010",
         713 => x"58010010",
         714 => x"58010010",
         715 => x"58010010",
         716 => x"58010010",
         717 => x"2c010010",
         718 => x"0d0a5448",
         719 => x"55415320",
         720 => x"52495343",
         721 => x"2d562042",
         722 => x"6f6f746c",
         723 => x"6f616465",
         724 => x"72207630",
         725 => x"2e322e31",
         726 => x"0d0a0000",
         727 => x"3f0a0000",
         728 => x"3e200000",
         729 => x"68000000",
         730 => x"48656c70",
         731 => x"3a0d0a20",
         732 => x"68202020",
         733 => x"20202020",
         734 => x"20202020",
         735 => x"20202020",
         736 => x"202d2074",
         737 => x"68697320",
         738 => x"68656c70",
         739 => x"0d0a2072",
         740 => x"20202020",
         741 => x"20202020",
         742 => x"20202020",
         743 => x"20202020",
         744 => x"2d207275",
         745 => x"6e206170",
         746 => x"706c6963",
         747 => x"6174696f",
         748 => x"6e0d0a20",
         749 => x"7277203c",
         750 => x"61646472",
         751 => x"3e202020",
         752 => x"20202020",
         753 => x"202d2072",
         754 => x"65616420",
         755 => x"776f7264",
         756 => x"2066726f",
         757 => x"6d206164",
         758 => x"64720d0a",
         759 => x"20777720",
         760 => x"3c616464",
         761 => x"723e203c",
         762 => x"64617461",
         763 => x"3e202d20",
         764 => x"77726974",
         765 => x"6520776f",
         766 => x"72642064",
         767 => x"61746120",
         768 => x"61742061",
         769 => x"6464720d",
         770 => x"0a206477",
         771 => x"203c6164",
         772 => x"64723e20",
         773 => x"20202020",
         774 => x"2020202d",
         775 => x"2064756d",
         776 => x"70203136",
         777 => x"20776f72",
         778 => x"64730d0a",
         779 => x"206e2020",
         780 => x"20202020",
         781 => x"20202020",
         782 => x"20202020",
         783 => x"20202d20",
         784 => x"64756d70",
         785 => x"206e6578",
         786 => x"74203136",
         787 => x"20776f72",
         788 => x"64730000",
         789 => x"72000000",
         790 => x"72772000",
         791 => x"3a200000",
         792 => x"4e6f7420",
         793 => x"6f6e2034",
         794 => x"2d627974",
         795 => x"6520626f",
         796 => x"756e6461",
         797 => x"72792100",
         798 => x"77772000",
         799 => x"64772000",
         800 => x"20200000",
         801 => x"3f3f0000",
         802 => x"626f6f74",
         803 => x"6c6f6164",
         804 => x"65720000",
         805 => x"54485541",
         806 => x"53205249",
         807 => x"53432d56",
         808 => x"20525633",
         809 => x"32494d20",
         810 => x"62617265",
         811 => x"206d6574",
         812 => x"616c2070",
         813 => x"726f6365",
         814 => x"73736f72",
         815 => x"00000000",
         816 => x"54686520",
         817 => x"48616775",
         818 => x"6520556e",
         819 => x"69766572",
         820 => x"73697479",
         821 => x"206f6620",
         822 => x"4170706c",
         823 => x"69656420",
         824 => x"53636965",
         825 => x"6e636573",
         826 => x"00000000",
         827 => x"44657061",
         828 => x"72746d65",
         829 => x"6e74206f",
         830 => x"6620456c",
         831 => x"65637472",
         832 => x"6963616c",
         833 => x"20456e67",
         834 => x"696e6565",
         835 => x"72696e67",
         836 => x"00000000",
         837 => x"4a2e452e",
         838 => x"4a2e206f",
         839 => x"70206465",
         840 => x"6e204272",
         841 => x"6f757700",
         842 => x"3c627265",
         843 => x"616b3e0d",
         844 => x"0a000000",
         845 => x"00202020",
         846 => x"20202020",
         847 => x"20202828",
         848 => x"28282820",
         849 => x"20202020",
         850 => x"20202020",
         851 => x"20202020",
         852 => x"20202020",
         853 => x"20881010",
         854 => x"10101010",
         855 => x"10101010",
         856 => x"10101010",
         857 => x"10040404",
         858 => x"04040404",
         859 => x"04040410",
         860 => x"10101010",
         861 => x"10104141",
         862 => x"41414141",
         863 => x"01010101",
         864 => x"01010101",
         865 => x"01010101",
         866 => x"01010101",
         867 => x"01010101",
         868 => x"10101010",
         869 => x"10104242",
         870 => x"42424242",
         871 => x"02020202",
         872 => x"02020202",
         873 => x"02020202",
         874 => x"02020202",
         875 => x"02020202",
         876 => x"10101010",
         877 => x"20000000",
         878 => x"00000000",
         879 => x"00000000",
         880 => x"00000000",
         881 => x"00000000",
         882 => x"00000000",
         883 => x"00000000",
         884 => x"00000000",
         885 => x"00000000",
         886 => x"00000000",
         887 => x"00000000",
         888 => x"00000000",
         889 => x"00000000",
         890 => x"00000000",
         891 => x"00000000",
         892 => x"00000000",
         893 => x"00000000",
         894 => x"00000000",
         895 => x"00000000",
         896 => x"00000000",
         897 => x"00000000",
         898 => x"00000000",
         899 => x"00000000",
         900 => x"00000000",
         901 => x"00000000",
         902 => x"00000000",
         903 => x"00000000",
         904 => x"00000000",
         905 => x"00000000",
         906 => x"00000000",
         907 => x"00000000",
         908 => x"00000000",
         909 => x"00000000",
         910 => x"18000020",
         911 => x"880c0010",
         912 => x"940c0010",
         913 => x"c00c0010",
         914 => x"ec0c0010",
         915 => x"140d0010",
         916 => x"00000000",
         917 => x"00000000",
         918 => x"00000000",
         919 => x"00000000",
         920 => x"00000000",
         921 => x"00000000",
         922 => x"00000000",
         923 => x"00000000",
         924 => x"00000000",
         925 => x"00000000",
         926 => x"00000000",
         927 => x"00000000",
         928 => x"00000000",
         929 => x"00000000",
         930 => x"00000000",
         931 => x"00000000",
         932 => x"00000000",
         933 => x"00000000",
         934 => x"00000000",
         935 => x"00000000",
         936 => x"00000000",
         937 => x"00000000",
         938 => x"00000000",
         939 => x"00000000",
         940 => x"00000000",
         941 => x"18000020",
         others => (others => '0')
        );

begin

    gen_bootrom: if HAVE_BOOTLOADER_ROM generate
        O_instruction_misaligned_error <= '0' when I_pc(1 downto 0) = "00" else '1';        

        -- ROM, for both instructions and read-only data
        process (I_clk, I_areset, I_pc, I_memaddress, I_csboot, I_memsize, I_stall) is
        variable address_instr : integer range 0 to bootloader_size-1;
        variable address_data : integer range 0 to bootloader_size-1;
        variable instr_var : data_type;
        variable instr_recode : data_type;
        variable romdata_var : data_type;
        constant x : data_type := (others => 'X');
        begin
            -- Calculate addresses
            address_instr := to_integer(unsigned(I_pc(bootloader_size_bits-1 downto 2)));
            address_data := to_integer(unsigned(I_memaddress(bootloader_size_bits-1 downto 2)));

            -- Quartus will detect ROM table and uses onboard RAM
            -- Do not use reset, otherwise ROM will be created with ALMs
            if rising_edge(I_clk) then
                if I_stall = '0' then
                    instr_var := bootrom(address_instr);
                end if;
                romdata_var := bootrom(address_data);
            end if;
            
            -- Recode instruction
            O_instr <= instr_var(7 downto 0) & instr_var(15 downto 8) & instr_var(23 downto 16) & instr_var(31 downto 24);
            
            O_load_misaligned_error <= '0';
            
            -- By natural size, for data
            if I_csboot = '1' then
                if I_memsize = memsize_word and I_memaddress(1 downto 0) = "00" then
                    O_dataout <= romdata_var(7 downto 0) & romdata_var(15 downto 8) & romdata_var(23 downto 16) & romdata_var(31 downto 24);
                elsif I_memsize = memsize_halfword and I_memaddress(1 downto 0) = "00" then
                    O_dataout <= x(31 downto 16) & romdata_var(23 downto 16) & romdata_var(31 downto 24);
                elsif I_memsize = memsize_halfword and I_memaddress(1 downto 0) = "10" then
                    O_dataout <= x(31 downto 16) & romdata_var(7 downto 0) & romdata_var(15 downto 8);
                elsif I_memsize = memsize_byte then
                    case I_memaddress(1 downto 0) is
                        when "00" => O_dataout <= x(31 downto 8) & romdata_var(31 downto 24);
                        when "01" => O_dataout <= x(31 downto 8) & romdata_var(23 downto 16);
                        when "10" => O_dataout <= x(31 downto 8) & romdata_var(15 downto 8);
                        when "11" => O_dataout <= x(31 downto 8) & romdata_var(7 downto 0);
                        when others => O_dataout <= x; O_load_misaligned_error <= '1';
                    end case;
                else
                    -- Chip select, but not aligned
                    O_dataout <= x;
                    O_load_misaligned_error <= '1';
                end if;
            else
                -- No chip select, so no data
                O_dataout <= x;
            end if;
        end process;
    end generate;

    gen_bootrom_not: if not HAVE_BOOTLOADER_ROM generate
        O_instruction_misaligned_error <= '0';
        O_load_misaligned_error <= '0';
        O_dataout <= (others => 'X');
        O_instr  <= (others => 'X');
    end generate;
end architecture rtl;
